library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;         --arquivo deve ser adicionado ao projeto

entity tabela_sin is
    generic (-- constant THETA_MAX : integer := 380808000;  --eqquivalente a 2*pi
                  constant n_bits_phase : integer :=16;  --numero de bits que representa a fase da rede
                  constant n_bits_c: integer := 16;  --numero de bits da portadora  
						constant I : integer := 1;  --número de bits da parte inteira excluindo sinal
						constant F : integer := 14 --número de bits da parte fracinária  
             );
   port(
		clk : in std_logic;
		theta: in std_logic_vector(15 downto 0);
		MAX :  in sfixed(15 downto 0); -- valor de contagem maximo 16 bits em sQ15.0
		ma : in sfixed(I downto -F); -- Indice de modulação em Q15
		va : out std_logic_vector(15 downto 0) -- Razão ciclica em Q0
	);
end tabela_sin;

architecture tabela_sin of tabela_sin is
    signal id : std_logic_vector(10 downto 0);
    signal sin : sfixed(I downto -F);
	 signal va_Q14 : sfixed(1 downto -14);  -- signed Q13
begin 
    
  id <= theta(n_bits_phase-1 downto n_bits_phase-11); -- 15 downto 5 - resolução do pwm?
   -- id <= theta; 
-- MAX == to_sfixed(1335,16,0);
	 
    process(clk)
    begin
        if rising_edge(clk) then		  
				va_Q14 <= resize((resize(sin*ma, 1, -14)+ to_sfixed(1, 1, -14)),1,-14); -- Valor entre +-1
				va <= to_slv(resize(va_Q14*scalb(MAX, -1),15,0)); --			
        end if;
    end process;
with id select
  sin <=  to_sfixed(0.000000,  I, -F) when "00000000000", 
		    to_sfixed(0.003068,  I, -F) when "00000000001", 
		    to_sfixed(0.006136,  I, -F) when "00000000010", 
		    to_sfixed(0.009204,  I, -F) when "00000000011", 
		    to_sfixed(0.012272,  I, -F) when "00000000100", 
		    to_sfixed(0.015339,  I, -F) when "00000000101", 
		    to_sfixed(0.018407,  I, -F) when "00000000110", 
		    to_sfixed(0.021474,  I, -F) when "00000000111", 
		    to_sfixed(0.024541,  I, -F) when "00000001000", 
		    to_sfixed(0.027608,  I, -F) when "00000001001", 
		    to_sfixed(0.030675,  I, -F) when "00000001010", 
		    to_sfixed(0.033741,  I, -F) when "00000001011", 
		    to_sfixed(0.036807,  I, -F) when "00000001100", 
		    to_sfixed(0.039873,  I, -F) when "00000001101", 
		    to_sfixed(0.042938,  I, -F) when "00000001110", 
		    to_sfixed(0.046003,  I, -F) when "00000001111", 
		    to_sfixed(0.049068,  I, -F) when "00000010000", 
		    to_sfixed(0.052132,  I, -F) when "00000010001", 
		    to_sfixed(0.055195,  I, -F) when "00000010010", 
		    to_sfixed(0.058258,  I, -F) when "00000010011", 
		    to_sfixed(0.061321,  I, -F) when "00000010100", 
		    to_sfixed(0.064383,  I, -F) when "00000010101", 
		    to_sfixed(0.067444,  I, -F) when "00000010110", 
		    to_sfixed(0.070505,  I, -F) when "00000010111", 
		    to_sfixed(0.073565,  I, -F) when "00000011000", 
		    to_sfixed(0.076624,  I, -F) when "00000011001", 
		    to_sfixed(0.079682,  I, -F) when "00000011010", 
		    to_sfixed(0.082740,  I, -F) when "00000011011", 
		    to_sfixed(0.085797,  I, -F) when "00000011100", 
		    to_sfixed(0.088854,  I, -F) when "00000011101", 
		    to_sfixed(0.091909,  I, -F) when "00000011110", 
		    to_sfixed(0.094963,  I, -F) when "00000011111", 
		    to_sfixed(0.098017,  I, -F) when "00000100000", 
		    to_sfixed(0.101070,  I, -F) when "00000100001", 
		    to_sfixed(0.104122,  I, -F) when "00000100010", 
		    to_sfixed(0.107172,  I, -F) when "00000100011", 
		    to_sfixed(0.110222,  I, -F) when "00000100100", 
		    to_sfixed(0.113271,  I, -F) when "00000100101", 
		    to_sfixed(0.116319,  I, -F) when "00000100110", 
		    to_sfixed(0.119365,  I, -F) when "00000100111", 
		    to_sfixed(0.122411,  I, -F) when "00000101000", 
		    to_sfixed(0.125455,  I, -F) when "00000101001", 
		    to_sfixed(0.128498,  I, -F) when "00000101010", 
		    to_sfixed(0.131540,  I, -F) when "00000101011", 
		    to_sfixed(0.134581,  I, -F) when "00000101100", 
		    to_sfixed(0.137620,  I, -F) when "00000101101", 
		    to_sfixed(0.140658,  I, -F) when "00000101110", 
		    to_sfixed(0.143695,  I, -F) when "00000101111", 
		    to_sfixed(0.146730,  I, -F) when "00000110000", 
		    to_sfixed(0.149765,  I, -F) when "00000110001", 
		    to_sfixed(0.152797,  I, -F) when "00000110010", 
		    to_sfixed(0.155828,  I, -F) when "00000110011", 
		    to_sfixed(0.158858,  I, -F) when "00000110100", 
		    to_sfixed(0.161886,  I, -F) when "00000110101", 
		    to_sfixed(0.164913,  I, -F) when "00000110110", 
		    to_sfixed(0.167938,  I, -F) when "00000110111", 
		    to_sfixed(0.170962,  I, -F) when "00000111000", 
		    to_sfixed(0.173984,  I, -F) when "00000111001", 
		    to_sfixed(0.177004,  I, -F) when "00000111010", 
		    to_sfixed(0.180023,  I, -F) when "00000111011", 
		    to_sfixed(0.183040,  I, -F) when "00000111100", 
		    to_sfixed(0.186055,  I, -F) when "00000111101", 
		    to_sfixed(0.189069,  I, -F) when "00000111110", 
		    to_sfixed(0.192080,  I, -F) when "00000111111", 
		    to_sfixed(0.195090,  I, -F) when "00001000000", 
		    to_sfixed(0.198098,  I, -F) when "00001000001", 
		    to_sfixed(0.201105,  I, -F) when "00001000010", 
		    to_sfixed(0.204109,  I, -F) when "00001000011", 
		    to_sfixed(0.207111,  I, -F) when "00001000100", 
		    to_sfixed(0.210112,  I, -F) when "00001000101", 
		    to_sfixed(0.213110,  I, -F) when "00001000110", 
		    to_sfixed(0.216107,  I, -F) when "00001000111", 
		    to_sfixed(0.219101,  I, -F) when "00001001000", 
		    to_sfixed(0.222094,  I, -F) when "00001001001", 
		    to_sfixed(0.225084,  I, -F) when "00001001010", 
		    to_sfixed(0.228072,  I, -F) when "00001001011", 
		    to_sfixed(0.231058,  I, -F) when "00001001100", 
		    to_sfixed(0.234042,  I, -F) when "00001001101", 
		    to_sfixed(0.237024,  I, -F) when "00001001110", 
		    to_sfixed(0.240003,  I, -F) when "00001001111", 
		    to_sfixed(0.242980,  I, -F) when "00001010000", 
		    to_sfixed(0.245955,  I, -F) when "00001010001", 
		    to_sfixed(0.248928,  I, -F) when "00001010010", 
		    to_sfixed(0.251898,  I, -F) when "00001010011", 
		    to_sfixed(0.254866,  I, -F) when "00001010100", 
		    to_sfixed(0.257831,  I, -F) when "00001010101", 
		    to_sfixed(0.260794,  I, -F) when "00001010110", 
		    to_sfixed(0.263755,  I, -F) when "00001010111", 
		    to_sfixed(0.266713,  I, -F) when "00001011000", 
		    to_sfixed(0.269668,  I, -F) when "00001011001", 
		    to_sfixed(0.272621,  I, -F) when "00001011010", 
		    to_sfixed(0.275572,  I, -F) when "00001011011", 
		    to_sfixed(0.278520,  I, -F) when "00001011100", 
		    to_sfixed(0.281465,  I, -F) when "00001011101", 
		    to_sfixed(0.284408,  I, -F) when "00001011110", 
		    to_sfixed(0.287347,  I, -F) when "00001011111", 
		    to_sfixed(0.290285,  I, -F) when "00001100000", 
		    to_sfixed(0.293219,  I, -F) when "00001100001", 
		    to_sfixed(0.296151,  I, -F) when "00001100010", 
		    to_sfixed(0.299080,  I, -F) when "00001100011", 
		    to_sfixed(0.302006,  I, -F) when "00001100100", 
		    to_sfixed(0.304929,  I, -F) when "00001100101", 
		    to_sfixed(0.307850,  I, -F) when "00001100110", 
		    to_sfixed(0.310767,  I, -F) when "00001100111", 
		    to_sfixed(0.313682,  I, -F) when "00001101000", 
		    to_sfixed(0.316593,  I, -F) when "00001101001", 
		    to_sfixed(0.319502,  I, -F) when "00001101010", 
		    to_sfixed(0.322408,  I, -F) when "00001101011", 
		    to_sfixed(0.325310,  I, -F) when "00001101100", 
		    to_sfixed(0.328210,  I, -F) when "00001101101", 
		    to_sfixed(0.331106,  I, -F) when "00001101110", 
		    to_sfixed(0.334000,  I, -F) when "00001101111", 
		    to_sfixed(0.336890,  I, -F) when "00001110000", 
		    to_sfixed(0.339777,  I, -F) when "00001110001", 
		    to_sfixed(0.342661,  I, -F) when "00001110010", 
		    to_sfixed(0.345541,  I, -F) when "00001110011", 
		    to_sfixed(0.348419,  I, -F) when "00001110100", 
		    to_sfixed(0.351293,  I, -F) when "00001110101", 
		    to_sfixed(0.354164,  I, -F) when "00001110110", 
		    to_sfixed(0.357031,  I, -F) when "00001110111", 
		    to_sfixed(0.359895,  I, -F) when "00001111000", 
		    to_sfixed(0.362756,  I, -F) when "00001111001", 
		    to_sfixed(0.365613,  I, -F) when "00001111010", 
		    to_sfixed(0.368467,  I, -F) when "00001111011", 
		    to_sfixed(0.371317,  I, -F) when "00001111100", 
		    to_sfixed(0.374164,  I, -F) when "00001111101", 
		    to_sfixed(0.377007,  I, -F) when "00001111110", 
		    to_sfixed(0.379847,  I, -F) when "00001111111", 
		    to_sfixed(0.382683,  I, -F) when "00010000000", 
		    to_sfixed(0.385516,  I, -F) when "00010000001", 
		    to_sfixed(0.388345,  I, -F) when "00010000010", 
		    to_sfixed(0.391170,  I, -F) when "00010000011", 
		    to_sfixed(0.393992,  I, -F) when "00010000100", 
		    to_sfixed(0.396810,  I, -F) when "00010000101", 
		    to_sfixed(0.399624,  I, -F) when "00010000110", 
		    to_sfixed(0.402435,  I, -F) when "00010000111", 
		    to_sfixed(0.405241,  I, -F) when "00010001000", 
		    to_sfixed(0.408044,  I, -F) when "00010001001", 
		    to_sfixed(0.410843,  I, -F) when "00010001010", 
		    to_sfixed(0.413638,  I, -F) when "00010001011", 
		    to_sfixed(0.416430,  I, -F) when "00010001100", 
		    to_sfixed(0.419217,  I, -F) when "00010001101", 
		    to_sfixed(0.422000,  I, -F) when "00010001110", 
		    to_sfixed(0.424780,  I, -F) when "00010001111", 
		    to_sfixed(0.427555,  I, -F) when "00010010000", 
		    to_sfixed(0.430326,  I, -F) when "00010010001", 
		    to_sfixed(0.433094,  I, -F) when "00010010010", 
		    to_sfixed(0.435857,  I, -F) when "00010010011", 
		    to_sfixed(0.438616,  I, -F) when "00010010100", 
		    to_sfixed(0.441371,  I, -F) when "00010010101", 
		    to_sfixed(0.444122,  I, -F) when "00010010110", 
		    to_sfixed(0.446869,  I, -F) when "00010010111", 
		    to_sfixed(0.449611,  I, -F) when "00010011000", 
		    to_sfixed(0.452350,  I, -F) when "00010011001", 
		    to_sfixed(0.455084,  I, -F) when "00010011010", 
		    to_sfixed(0.457813,  I, -F) when "00010011011", 
		    to_sfixed(0.460539,  I, -F) when "00010011100", 
		    to_sfixed(0.463260,  I, -F) when "00010011101", 
		    to_sfixed(0.465976,  I, -F) when "00010011110", 
		    to_sfixed(0.468689,  I, -F) when "00010011111", 
		    to_sfixed(0.471397,  I, -F) when "00010100000", 
		    to_sfixed(0.474100,  I, -F) when "00010100001", 
		    to_sfixed(0.476799,  I, -F) when "00010100010", 
		    to_sfixed(0.479494,  I, -F) when "00010100011", 
		    to_sfixed(0.482184,  I, -F) when "00010100100", 
		    to_sfixed(0.484869,  I, -F) when "00010100101", 
		    to_sfixed(0.487550,  I, -F) when "00010100110", 
		    to_sfixed(0.490226,  I, -F) when "00010100111", 
		    to_sfixed(0.492898,  I, -F) when "00010101000", 
		    to_sfixed(0.495565,  I, -F) when "00010101001", 
		    to_sfixed(0.498228,  I, -F) when "00010101010", 
		    to_sfixed(0.500885,  I, -F) when "00010101011", 
		    to_sfixed(0.503538,  I, -F) when "00010101100", 
		    to_sfixed(0.506187,  I, -F) when "00010101101", 
		    to_sfixed(0.508830,  I, -F) when "00010101110", 
		    to_sfixed(0.511469,  I, -F) when "00010101111", 
		    to_sfixed(0.514103,  I, -F) when "00010110000", 
		    to_sfixed(0.516732,  I, -F) when "00010110001", 
		    to_sfixed(0.519356,  I, -F) when "00010110010", 
		    to_sfixed(0.521975,  I, -F) when "00010110011", 
		    to_sfixed(0.524590,  I, -F) when "00010110100", 
		    to_sfixed(0.527199,  I, -F) when "00010110101", 
		    to_sfixed(0.529804,  I, -F) when "00010110110", 
		    to_sfixed(0.532403,  I, -F) when "00010110111", 
		    to_sfixed(0.534998,  I, -F) when "00010111000", 
		    to_sfixed(0.537587,  I, -F) when "00010111001", 
		    to_sfixed(0.540171,  I, -F) when "00010111010", 
		    to_sfixed(0.542751,  I, -F) when "00010111011", 
		    to_sfixed(0.545325,  I, -F) when "00010111100", 
		    to_sfixed(0.547894,  I, -F) when "00010111101", 
		    to_sfixed(0.550458,  I, -F) when "00010111110", 
		    to_sfixed(0.553017,  I, -F) when "00010111111", 
		    to_sfixed(0.555570,  I, -F) when "00011000000", 
		    to_sfixed(0.558119,  I, -F) when "00011000001", 
		    to_sfixed(0.560662,  I, -F) when "00011000010", 
		    to_sfixed(0.563199,  I, -F) when "00011000011", 
		    to_sfixed(0.565732,  I, -F) when "00011000100", 
		    to_sfixed(0.568259,  I, -F) when "00011000101", 
		    to_sfixed(0.570781,  I, -F) when "00011000110", 
		    to_sfixed(0.573297,  I, -F) when "00011000111", 
		    to_sfixed(0.575808,  I, -F) when "00011001000", 
		    to_sfixed(0.578314,  I, -F) when "00011001001", 
		    to_sfixed(0.580814,  I, -F) when "00011001010", 
		    to_sfixed(0.583309,  I, -F) when "00011001011", 
		    to_sfixed(0.585798,  I, -F) when "00011001100", 
		    to_sfixed(0.588282,  I, -F) when "00011001101", 
		    to_sfixed(0.590760,  I, -F) when "00011001110", 
		    to_sfixed(0.593232,  I, -F) when "00011001111", 
		    to_sfixed(0.595699,  I, -F) when "00011010000", 
		    to_sfixed(0.598161,  I, -F) when "00011010001", 
		    to_sfixed(0.600616,  I, -F) when "00011010010", 
		    to_sfixed(0.603067,  I, -F) when "00011010011", 
		    to_sfixed(0.605511,  I, -F) when "00011010100", 
		    to_sfixed(0.607950,  I, -F) when "00011010101", 
		    to_sfixed(0.610383,  I, -F) when "00011010110", 
		    to_sfixed(0.612810,  I, -F) when "00011010111", 
		    to_sfixed(0.615232,  I, -F) when "00011011000", 
		    to_sfixed(0.617647,  I, -F) when "00011011001", 
		    to_sfixed(0.620057,  I, -F) when "00011011010", 
		    to_sfixed(0.622461,  I, -F) when "00011011011", 
		    to_sfixed(0.624859,  I, -F) when "00011011100", 
		    to_sfixed(0.627252,  I, -F) when "00011011101", 
		    to_sfixed(0.629638,  I, -F) when "00011011110", 
		    to_sfixed(0.632019,  I, -F) when "00011011111", 
		    to_sfixed(0.634393,  I, -F) when "00011100000", 
		    to_sfixed(0.636762,  I, -F) when "00011100001", 
		    to_sfixed(0.639124,  I, -F) when "00011100010", 
		    to_sfixed(0.641481,  I, -F) when "00011100011", 
		    to_sfixed(0.643832,  I, -F) when "00011100100", 
		    to_sfixed(0.646176,  I, -F) when "00011100101", 
		    to_sfixed(0.648514,  I, -F) when "00011100110", 
		    to_sfixed(0.650847,  I, -F) when "00011100111", 
		    to_sfixed(0.653173,  I, -F) when "00011101000", 
		    to_sfixed(0.655493,  I, -F) when "00011101001", 
		    to_sfixed(0.657807,  I, -F) when "00011101010", 
		    to_sfixed(0.660114,  I, -F) when "00011101011", 
		    to_sfixed(0.662416,  I, -F) when "00011101100", 
		    to_sfixed(0.664711,  I, -F) when "00011101101", 
		    to_sfixed(0.667000,  I, -F) when "00011101110", 
		    to_sfixed(0.669283,  I, -F) when "00011101111", 
		    to_sfixed(0.671559,  I, -F) when "00011110000", 
		    to_sfixed(0.673829,  I, -F) when "00011110001", 
		    to_sfixed(0.676093,  I, -F) when "00011110010", 
		    to_sfixed(0.678350,  I, -F) when "00011110011", 
		    to_sfixed(0.680601,  I, -F) when "00011110100", 
		    to_sfixed(0.682846,  I, -F) when "00011110101", 
		    to_sfixed(0.685084,  I, -F) when "00011110110", 
		    to_sfixed(0.687315,  I, -F) when "00011110111", 
		    to_sfixed(0.689541,  I, -F) when "00011111000", 
		    to_sfixed(0.691759,  I, -F) when "00011111001", 
		    to_sfixed(0.693971,  I, -F) when "00011111010", 
		    to_sfixed(0.696177,  I, -F) when "00011111011", 
		    to_sfixed(0.698376,  I, -F) when "00011111100", 
		    to_sfixed(0.700569,  I, -F) when "00011111101", 
		    to_sfixed(0.702755,  I, -F) when "00011111110", 
		    to_sfixed(0.704934,  I, -F) when "00011111111", 
		    to_sfixed(0.707107,  I, -F) when "00100000000", 
		    to_sfixed(0.709273,  I, -F) when "00100000001", 
		    to_sfixed(0.711432,  I, -F) when "00100000010", 
		    to_sfixed(0.713585,  I, -F) when "00100000011", 
		    to_sfixed(0.715731,  I, -F) when "00100000100", 
		    to_sfixed(0.717870,  I, -F) when "00100000101", 
		    to_sfixed(0.720003,  I, -F) when "00100000110", 
		    to_sfixed(0.722128,  I, -F) when "00100000111", 
		    to_sfixed(0.724247,  I, -F) when "00100001000", 
		    to_sfixed(0.726359,  I, -F) when "00100001001", 
		    to_sfixed(0.728464,  I, -F) when "00100001010", 
		    to_sfixed(0.730563,  I, -F) when "00100001011", 
		    to_sfixed(0.732654,  I, -F) when "00100001100", 
		    to_sfixed(0.734739,  I, -F) when "00100001101", 
		    to_sfixed(0.736817,  I, -F) when "00100001110", 
		    to_sfixed(0.738887,  I, -F) when "00100001111", 
		    to_sfixed(0.740951,  I, -F) when "00100010000", 
		    to_sfixed(0.743008,  I, -F) when "00100010001", 
		    to_sfixed(0.745058,  I, -F) when "00100010010", 
		    to_sfixed(0.747101,  I, -F) when "00100010011", 
		    to_sfixed(0.749136,  I, -F) when "00100010100", 
		    to_sfixed(0.751165,  I, -F) when "00100010101", 
		    to_sfixed(0.753187,  I, -F) when "00100010110", 
		    to_sfixed(0.755201,  I, -F) when "00100010111", 
		    to_sfixed(0.757209,  I, -F) when "00100011000", 
		    to_sfixed(0.759209,  I, -F) when "00100011001", 
		    to_sfixed(0.761202,  I, -F) when "00100011010", 
		    to_sfixed(0.763188,  I, -F) when "00100011011", 
		    to_sfixed(0.765167,  I, -F) when "00100011100", 
		    to_sfixed(0.767139,  I, -F) when "00100011101", 
		    to_sfixed(0.769103,  I, -F) when "00100011110", 
		    to_sfixed(0.771061,  I, -F) when "00100011111", 
		    to_sfixed(0.773010,  I, -F) when "00100100000", 
		    to_sfixed(0.774953,  I, -F) when "00100100001", 
		    to_sfixed(0.776888,  I, -F) when "00100100010", 
		    to_sfixed(0.778817,  I, -F) when "00100100011", 
		    to_sfixed(0.780737,  I, -F) when "00100100100", 
		    to_sfixed(0.782651,  I, -F) when "00100100101", 
		    to_sfixed(0.784557,  I, -F) when "00100100110", 
		    to_sfixed(0.786455,  I, -F) when "00100100111", 
		    to_sfixed(0.788346,  I, -F) when "00100101000", 
		    to_sfixed(0.790230,  I, -F) when "00100101001", 
		    to_sfixed(0.792107,  I, -F) when "00100101010", 
		    to_sfixed(0.793975,  I, -F) when "00100101011", 
		    to_sfixed(0.795837,  I, -F) when "00100101100", 
		    to_sfixed(0.797691,  I, -F) when "00100101101", 
		    to_sfixed(0.799537,  I, -F) when "00100101110", 
		    to_sfixed(0.801376,  I, -F) when "00100101111", 
		    to_sfixed(0.803208,  I, -F) when "00100110000", 
		    to_sfixed(0.805031,  I, -F) when "00100110001", 
		    to_sfixed(0.806848,  I, -F) when "00100110010", 
		    to_sfixed(0.808656,  I, -F) when "00100110011", 
		    to_sfixed(0.810457,  I, -F) when "00100110100", 
		    to_sfixed(0.812251,  I, -F) when "00100110101", 
		    to_sfixed(0.814036,  I, -F) when "00100110110", 
		    to_sfixed(0.815814,  I, -F) when "00100110111", 
		    to_sfixed(0.817585,  I, -F) when "00100111000", 
		    to_sfixed(0.819348,  I, -F) when "00100111001", 
		    to_sfixed(0.821103,  I, -F) when "00100111010", 
		    to_sfixed(0.822850,  I, -F) when "00100111011", 
		    to_sfixed(0.824589,  I, -F) when "00100111100", 
		    to_sfixed(0.826321,  I, -F) when "00100111101", 
		    to_sfixed(0.828045,  I, -F) when "00100111110", 
		    to_sfixed(0.829761,  I, -F) when "00100111111", 
		    to_sfixed(0.831470,  I, -F) when "00101000000", 
		    to_sfixed(0.833170,  I, -F) when "00101000001", 
		    to_sfixed(0.834863,  I, -F) when "00101000010", 
		    to_sfixed(0.836548,  I, -F) when "00101000011", 
		    to_sfixed(0.838225,  I, -F) when "00101000100", 
		    to_sfixed(0.839894,  I, -F) when "00101000101", 
		    to_sfixed(0.841555,  I, -F) when "00101000110", 
		    to_sfixed(0.843208,  I, -F) when "00101000111", 
		    to_sfixed(0.844854,  I, -F) when "00101001000", 
		    to_sfixed(0.846491,  I, -F) when "00101001001", 
		    to_sfixed(0.848120,  I, -F) when "00101001010", 
		    to_sfixed(0.849742,  I, -F) when "00101001011", 
		    to_sfixed(0.851355,  I, -F) when "00101001100", 
		    to_sfixed(0.852961,  I, -F) when "00101001101", 
		    to_sfixed(0.854558,  I, -F) when "00101001110", 
		    to_sfixed(0.856147,  I, -F) when "00101001111", 
		    to_sfixed(0.857729,  I, -F) when "00101010000", 
		    to_sfixed(0.859302,  I, -F) when "00101010001", 
		    to_sfixed(0.860867,  I, -F) when "00101010010", 
		    to_sfixed(0.862424,  I, -F) when "00101010011", 
		    to_sfixed(0.863973,  I, -F) when "00101010100", 
		    to_sfixed(0.865514,  I, -F) when "00101010101", 
		    to_sfixed(0.867046,  I, -F) when "00101010110", 
		    to_sfixed(0.868571,  I, -F) when "00101010111", 
		    to_sfixed(0.870087,  I, -F) when "00101011000", 
		    to_sfixed(0.871595,  I, -F) when "00101011001", 
		    to_sfixed(0.873095,  I, -F) when "00101011010", 
		    to_sfixed(0.874587,  I, -F) when "00101011011", 
		    to_sfixed(0.876070,  I, -F) when "00101011100", 
		    to_sfixed(0.877545,  I, -F) when "00101011101", 
		    to_sfixed(0.879012,  I, -F) when "00101011110", 
		    to_sfixed(0.880471,  I, -F) when "00101011111", 
		    to_sfixed(0.881921,  I, -F) when "00101100000", 
		    to_sfixed(0.883363,  I, -F) when "00101100001", 
		    to_sfixed(0.884797,  I, -F) when "00101100010", 
		    to_sfixed(0.886223,  I, -F) when "00101100011", 
		    to_sfixed(0.887640,  I, -F) when "00101100100", 
		    to_sfixed(0.889048,  I, -F) when "00101100101", 
		    to_sfixed(0.890449,  I, -F) when "00101100110", 
		    to_sfixed(0.891841,  I, -F) when "00101100111", 
		    to_sfixed(0.893224,  I, -F) when "00101101000", 
		    to_sfixed(0.894599,  I, -F) when "00101101001", 
		    to_sfixed(0.895966,  I, -F) when "00101101010", 
		    to_sfixed(0.897325,  I, -F) when "00101101011", 
		    to_sfixed(0.898674,  I, -F) when "00101101100", 
		    to_sfixed(0.900016,  I, -F) when "00101101101", 
		    to_sfixed(0.901349,  I, -F) when "00101101110", 
		    to_sfixed(0.902673,  I, -F) when "00101101111", 
		    to_sfixed(0.903989,  I, -F) when "00101110000", 
		    to_sfixed(0.905297,  I, -F) when "00101110001", 
		    to_sfixed(0.906596,  I, -F) when "00101110010", 
		    to_sfixed(0.907886,  I, -F) when "00101110011", 
		    to_sfixed(0.909168,  I, -F) when "00101110100", 
		    to_sfixed(0.910441,  I, -F) when "00101110101", 
		    to_sfixed(0.911706,  I, -F) when "00101110110", 
		    to_sfixed(0.912962,  I, -F) when "00101110111", 
		    to_sfixed(0.914210,  I, -F) when "00101111000", 
		    to_sfixed(0.915449,  I, -F) when "00101111001", 
		    to_sfixed(0.916679,  I, -F) when "00101111010", 
		    to_sfixed(0.917901,  I, -F) when "00101111011", 
		    to_sfixed(0.919114,  I, -F) when "00101111100", 
		    to_sfixed(0.920318,  I, -F) when "00101111101", 
		    to_sfixed(0.921514,  I, -F) when "00101111110", 
		    to_sfixed(0.922701,  I, -F) when "00101111111", 
		    to_sfixed(0.923880,  I, -F) when "00110000000", 
		    to_sfixed(0.925049,  I, -F) when "00110000001", 
		    to_sfixed(0.926210,  I, -F) when "00110000010", 
		    to_sfixed(0.927363,  I, -F) when "00110000011", 
		    to_sfixed(0.928506,  I, -F) when "00110000100", 
		    to_sfixed(0.929641,  I, -F) when "00110000101", 
		    to_sfixed(0.930767,  I, -F) when "00110000110", 
		    to_sfixed(0.931884,  I, -F) when "00110000111", 
		    to_sfixed(0.932993,  I, -F) when "00110001000", 
		    to_sfixed(0.934093,  I, -F) when "00110001001", 
		    to_sfixed(0.935184,  I, -F) when "00110001010", 
		    to_sfixed(0.936266,  I, -F) when "00110001011", 
		    to_sfixed(0.937339,  I, -F) when "00110001100", 
		    to_sfixed(0.938404,  I, -F) when "00110001101", 
		    to_sfixed(0.939459,  I, -F) when "00110001110", 
		    to_sfixed(0.940506,  I, -F) when "00110001111", 
		    to_sfixed(0.941544,  I, -F) when "00110010000", 
		    to_sfixed(0.942573,  I, -F) when "00110010001", 
		    to_sfixed(0.943593,  I, -F) when "00110010010", 
		    to_sfixed(0.944605,  I, -F) when "00110010011", 
		    to_sfixed(0.945607,  I, -F) when "00110010100", 
		    to_sfixed(0.946601,  I, -F) when "00110010101", 
		    to_sfixed(0.947586,  I, -F) when "00110010110", 
		    to_sfixed(0.948561,  I, -F) when "00110010111", 
		    to_sfixed(0.949528,  I, -F) when "00110011000", 
		    to_sfixed(0.950486,  I, -F) when "00110011001", 
		    to_sfixed(0.951435,  I, -F) when "00110011010", 
		    to_sfixed(0.952375,  I, -F) when "00110011011", 
		    to_sfixed(0.953306,  I, -F) when "00110011100", 
		    to_sfixed(0.954228,  I, -F) when "00110011101", 
		    to_sfixed(0.955141,  I, -F) when "00110011110", 
		    to_sfixed(0.956045,  I, -F) when "00110011111", 
		    to_sfixed(0.956940,  I, -F) when "00110100000", 
		    to_sfixed(0.957826,  I, -F) when "00110100001", 
		    to_sfixed(0.958703,  I, -F) when "00110100010", 
		    to_sfixed(0.959572,  I, -F) when "00110100011", 
		    to_sfixed(0.960431,  I, -F) when "00110100100", 
		    to_sfixed(0.961280,  I, -F) when "00110100101", 
		    to_sfixed(0.962121,  I, -F) when "00110100110", 
		    to_sfixed(0.962953,  I, -F) when "00110100111", 
		    to_sfixed(0.963776,  I, -F) when "00110101000", 
		    to_sfixed(0.964590,  I, -F) when "00110101001", 
		    to_sfixed(0.965394,  I, -F) when "00110101010", 
		    to_sfixed(0.966190,  I, -F) when "00110101011", 
		    to_sfixed(0.966976,  I, -F) when "00110101100", 
		    to_sfixed(0.967754,  I, -F) when "00110101101", 
		    to_sfixed(0.968522,  I, -F) when "00110101110", 
		    to_sfixed(0.969281,  I, -F) when "00110101111", 
		    to_sfixed(0.970031,  I, -F) when "00110110000", 
		    to_sfixed(0.970772,  I, -F) when "00110110001", 
		    to_sfixed(0.971504,  I, -F) when "00110110010", 
		    to_sfixed(0.972226,  I, -F) when "00110110011", 
		    to_sfixed(0.972940,  I, -F) when "00110110100", 
		    to_sfixed(0.973644,  I, -F) when "00110110101", 
		    to_sfixed(0.974339,  I, -F) when "00110110110", 
		    to_sfixed(0.975025,  I, -F) when "00110110111", 
		    to_sfixed(0.975702,  I, -F) when "00110111000", 
		    to_sfixed(0.976370,  I, -F) when "00110111001", 
		    to_sfixed(0.977028,  I, -F) when "00110111010", 
		    to_sfixed(0.977677,  I, -F) when "00110111011", 
		    to_sfixed(0.978317,  I, -F) when "00110111100", 
		    to_sfixed(0.978948,  I, -F) when "00110111101", 
		    to_sfixed(0.979570,  I, -F) when "00110111110", 
		    to_sfixed(0.980182,  I, -F) when "00110111111", 
		    to_sfixed(0.980785,  I, -F) when "00111000000", 
		    to_sfixed(0.981379,  I, -F) when "00111000001", 
		    to_sfixed(0.981964,  I, -F) when "00111000010", 
		    to_sfixed(0.982539,  I, -F) when "00111000011", 
		    to_sfixed(0.983105,  I, -F) when "00111000100", 
		    to_sfixed(0.983662,  I, -F) when "00111000101", 
		    to_sfixed(0.984210,  I, -F) when "00111000110", 
		    to_sfixed(0.984749,  I, -F) when "00111000111", 
		    to_sfixed(0.985278,  I, -F) when "00111001000", 
		    to_sfixed(0.985798,  I, -F) when "00111001001", 
		    to_sfixed(0.986308,  I, -F) when "00111001010", 
		    to_sfixed(0.986809,  I, -F) when "00111001011", 
		    to_sfixed(0.987301,  I, -F) when "00111001100", 
		    to_sfixed(0.987784,  I, -F) when "00111001101", 
		    to_sfixed(0.988258,  I, -F) when "00111001110", 
		    to_sfixed(0.988722,  I, -F) when "00111001111", 
		    to_sfixed(0.989177,  I, -F) when "00111010000", 
		    to_sfixed(0.989622,  I, -F) when "00111010001", 
		    to_sfixed(0.990058,  I, -F) when "00111010010", 
		    to_sfixed(0.990485,  I, -F) when "00111010011", 
		    to_sfixed(0.990903,  I, -F) when "00111010100", 
		    to_sfixed(0.991311,  I, -F) when "00111010101", 
		    to_sfixed(0.991710,  I, -F) when "00111010110", 
		    to_sfixed(0.992099,  I, -F) when "00111010111", 
		    to_sfixed(0.992480,  I, -F) when "00111011000", 
		    to_sfixed(0.992850,  I, -F) when "00111011001", 
		    to_sfixed(0.993212,  I, -F) when "00111011010", 
		    to_sfixed(0.993564,  I, -F) when "00111011011", 
		    to_sfixed(0.993907,  I, -F) when "00111011100", 
		    to_sfixed(0.994240,  I, -F) when "00111011101", 
		    to_sfixed(0.994565,  I, -F) when "00111011110", 
		    to_sfixed(0.994879,  I, -F) when "00111011111", 
		    to_sfixed(0.995185,  I, -F) when "00111100000", 
		    to_sfixed(0.995481,  I, -F) when "00111100001", 
		    to_sfixed(0.995767,  I, -F) when "00111100010", 
		    to_sfixed(0.996045,  I, -F) when "00111100011", 
		    to_sfixed(0.996313,  I, -F) when "00111100100", 
		    to_sfixed(0.996571,  I, -F) when "00111100101", 
		    to_sfixed(0.996820,  I, -F) when "00111100110", 
		    to_sfixed(0.997060,  I, -F) when "00111100111", 
		    to_sfixed(0.997290,  I, -F) when "00111101000", 
		    to_sfixed(0.997511,  I, -F) when "00111101001", 
		    to_sfixed(0.997723,  I, -F) when "00111101010", 
		    to_sfixed(0.997925,  I, -F) when "00111101011", 
		    to_sfixed(0.998118,  I, -F) when "00111101100", 
		    to_sfixed(0.998302,  I, -F) when "00111101101", 
		    to_sfixed(0.998476,  I, -F) when "00111101110", 
		    to_sfixed(0.998640,  I, -F) when "00111101111", 
		    to_sfixed(0.998795,  I, -F) when "00111110000", 
		    to_sfixed(0.998941,  I, -F) when "00111110001", 
		    to_sfixed(0.999078,  I, -F) when "00111110010", 
		    to_sfixed(0.999205,  I, -F) when "00111110011", 
		    to_sfixed(0.999322,  I, -F) when "00111110100", 
		    to_sfixed(0.999431,  I, -F) when "00111110101", 
		    to_sfixed(0.999529,  I, -F) when "00111110110", 
		    to_sfixed(0.999619,  I, -F) when "00111110111", 
		    to_sfixed(0.999699,  I, -F) when "00111111000", 
		    to_sfixed(0.999769,  I, -F) when "00111111001", 
		    to_sfixed(0.999831,  I, -F) when "00111111010", 
		    to_sfixed(0.999882,  I, -F) when "00111111011", 
		    to_sfixed(0.999925,  I, -F) when "00111111100", 
		    to_sfixed(0.999958,  I, -F) when "00111111101", 
		    to_sfixed(0.999981,  I, -F) when "00111111110", 
		    to_sfixed(0.999995,  I, -F) when "00111111111", 
		    to_sfixed(1.000000,  I, -F) when "01000000000", 
		    to_sfixed(0.999995,  I, -F) when "01000000001", 
		    to_sfixed(0.999981,  I, -F) when "01000000010", 
		    to_sfixed(0.999958,  I, -F) when "01000000011", 
		    to_sfixed(0.999925,  I, -F) when "01000000100", 
		    to_sfixed(0.999882,  I, -F) when "01000000101", 
		    to_sfixed(0.999831,  I, -F) when "01000000110", 
		    to_sfixed(0.999769,  I, -F) when "01000000111", 
		    to_sfixed(0.999699,  I, -F) when "01000001000", 
		    to_sfixed(0.999619,  I, -F) when "01000001001", 
		    to_sfixed(0.999529,  I, -F) when "01000001010", 
		    to_sfixed(0.999431,  I, -F) when "01000001011", 
		    to_sfixed(0.999322,  I, -F) when "01000001100", 
		    to_sfixed(0.999205,  I, -F) when "01000001101", 
		    to_sfixed(0.999078,  I, -F) when "01000001110", 
		    to_sfixed(0.998941,  I, -F) when "01000001111", 
		    to_sfixed(0.998795,  I, -F) when "01000010000", 
		    to_sfixed(0.998640,  I, -F) when "01000010001", 
		    to_sfixed(0.998476,  I, -F) when "01000010010", 
		    to_sfixed(0.998302,  I, -F) when "01000010011", 
		    to_sfixed(0.998118,  I, -F) when "01000010100", 
		    to_sfixed(0.997925,  I, -F) when "01000010101", 
		    to_sfixed(0.997723,  I, -F) when "01000010110", 
		    to_sfixed(0.997511,  I, -F) when "01000010111", 
		    to_sfixed(0.997290,  I, -F) when "01000011000", 
		    to_sfixed(0.997060,  I, -F) when "01000011001", 
		    to_sfixed(0.996820,  I, -F) when "01000011010", 
		    to_sfixed(0.996571,  I, -F) when "01000011011", 
		    to_sfixed(0.996313,  I, -F) when "01000011100", 
		    to_sfixed(0.996045,  I, -F) when "01000011101", 
		    to_sfixed(0.995767,  I, -F) when "01000011110", 
		    to_sfixed(0.995481,  I, -F) when "01000011111", 
		    to_sfixed(0.995185,  I, -F) when "01000100000", 
		    to_sfixed(0.994879,  I, -F) when "01000100001", 
		    to_sfixed(0.994565,  I, -F) when "01000100010", 
		    to_sfixed(0.994240,  I, -F) when "01000100011", 
		    to_sfixed(0.993907,  I, -F) when "01000100100", 
		    to_sfixed(0.993564,  I, -F) when "01000100101", 
		    to_sfixed(0.993212,  I, -F) when "01000100110", 
		    to_sfixed(0.992850,  I, -F) when "01000100111", 
		    to_sfixed(0.992480,  I, -F) when "01000101000", 
		    to_sfixed(0.992099,  I, -F) when "01000101001", 
		    to_sfixed(0.991710,  I, -F) when "01000101010", 
		    to_sfixed(0.991311,  I, -F) when "01000101011", 
		    to_sfixed(0.990903,  I, -F) when "01000101100", 
		    to_sfixed(0.990485,  I, -F) when "01000101101", 
		    to_sfixed(0.990058,  I, -F) when "01000101110", 
		    to_sfixed(0.989622,  I, -F) when "01000101111", 
		    to_sfixed(0.989177,  I, -F) when "01000110000", 
		    to_sfixed(0.988722,  I, -F) when "01000110001", 
		    to_sfixed(0.988258,  I, -F) when "01000110010", 
		    to_sfixed(0.987784,  I, -F) when "01000110011", 
		    to_sfixed(0.987301,  I, -F) when "01000110100", 
		    to_sfixed(0.986809,  I, -F) when "01000110101", 
		    to_sfixed(0.986308,  I, -F) when "01000110110", 
		    to_sfixed(0.985798,  I, -F) when "01000110111", 
		    to_sfixed(0.985278,  I, -F) when "01000111000", 
		    to_sfixed(0.984749,  I, -F) when "01000111001", 
		    to_sfixed(0.984210,  I, -F) when "01000111010", 
		    to_sfixed(0.983662,  I, -F) when "01000111011", 
		    to_sfixed(0.983105,  I, -F) when "01000111100", 
		    to_sfixed(0.982539,  I, -F) when "01000111101", 
		    to_sfixed(0.981964,  I, -F) when "01000111110", 
		    to_sfixed(0.981379,  I, -F) when "01000111111", 
		    to_sfixed(0.980785,  I, -F) when "01001000000", 
		    to_sfixed(0.980182,  I, -F) when "01001000001", 
		    to_sfixed(0.979570,  I, -F) when "01001000010", 
		    to_sfixed(0.978948,  I, -F) when "01001000011", 
		    to_sfixed(0.978317,  I, -F) when "01001000100", 
		    to_sfixed(0.977677,  I, -F) when "01001000101", 
		    to_sfixed(0.977028,  I, -F) when "01001000110", 
		    to_sfixed(0.976370,  I, -F) when "01001000111", 
		    to_sfixed(0.975702,  I, -F) when "01001001000", 
		    to_sfixed(0.975025,  I, -F) when "01001001001", 
		    to_sfixed(0.974339,  I, -F) when "01001001010", 
		    to_sfixed(0.973644,  I, -F) when "01001001011", 
		    to_sfixed(0.972940,  I, -F) when "01001001100", 
		    to_sfixed(0.972226,  I, -F) when "01001001101", 
		    to_sfixed(0.971504,  I, -F) when "01001001110", 
		    to_sfixed(0.970772,  I, -F) when "01001001111", 
		    to_sfixed(0.970031,  I, -F) when "01001010000", 
		    to_sfixed(0.969281,  I, -F) when "01001010001", 
		    to_sfixed(0.968522,  I, -F) when "01001010010", 
		    to_sfixed(0.967754,  I, -F) when "01001010011", 
		    to_sfixed(0.966976,  I, -F) when "01001010100", 
		    to_sfixed(0.966190,  I, -F) when "01001010101", 
		    to_sfixed(0.965394,  I, -F) when "01001010110", 
		    to_sfixed(0.964590,  I, -F) when "01001010111", 
		    to_sfixed(0.963776,  I, -F) when "01001011000", 
		    to_sfixed(0.962953,  I, -F) when "01001011001", 
		    to_sfixed(0.962121,  I, -F) when "01001011010", 
		    to_sfixed(0.961280,  I, -F) when "01001011011", 
		    to_sfixed(0.960431,  I, -F) when "01001011100", 
		    to_sfixed(0.959572,  I, -F) when "01001011101", 
		    to_sfixed(0.958703,  I, -F) when "01001011110", 
		    to_sfixed(0.957826,  I, -F) when "01001011111", 
		    to_sfixed(0.956940,  I, -F) when "01001100000", 
		    to_sfixed(0.956045,  I, -F) when "01001100001", 
		    to_sfixed(0.955141,  I, -F) when "01001100010", 
		    to_sfixed(0.954228,  I, -F) when "01001100011", 
		    to_sfixed(0.953306,  I, -F) when "01001100100", 
		    to_sfixed(0.952375,  I, -F) when "01001100101", 
		    to_sfixed(0.951435,  I, -F) when "01001100110", 
		    to_sfixed(0.950486,  I, -F) when "01001100111", 
		    to_sfixed(0.949528,  I, -F) when "01001101000", 
		    to_sfixed(0.948561,  I, -F) when "01001101001", 
		    to_sfixed(0.947586,  I, -F) when "01001101010", 
		    to_sfixed(0.946601,  I, -F) when "01001101011", 
		    to_sfixed(0.945607,  I, -F) when "01001101100", 
		    to_sfixed(0.944605,  I, -F) when "01001101101", 
		    to_sfixed(0.943593,  I, -F) when "01001101110", 
		    to_sfixed(0.942573,  I, -F) when "01001101111", 
		    to_sfixed(0.941544,  I, -F) when "01001110000", 
		    to_sfixed(0.940506,  I, -F) when "01001110001", 
		    to_sfixed(0.939459,  I, -F) when "01001110010", 
		    to_sfixed(0.938404,  I, -F) when "01001110011", 
		    to_sfixed(0.937339,  I, -F) when "01001110100", 
		    to_sfixed(0.936266,  I, -F) when "01001110101", 
		    to_sfixed(0.935184,  I, -F) when "01001110110", 
		    to_sfixed(0.934093,  I, -F) when "01001110111", 
		    to_sfixed(0.932993,  I, -F) when "01001111000", 
		    to_sfixed(0.931884,  I, -F) when "01001111001", 
		    to_sfixed(0.930767,  I, -F) when "01001111010", 
		    to_sfixed(0.929641,  I, -F) when "01001111011", 
		    to_sfixed(0.928506,  I, -F) when "01001111100", 
		    to_sfixed(0.927363,  I, -F) when "01001111101", 
		    to_sfixed(0.926210,  I, -F) when "01001111110", 
		    to_sfixed(0.925049,  I, -F) when "01001111111", 
		    to_sfixed(0.923880,  I, -F) when "01010000000", 
		    to_sfixed(0.922701,  I, -F) when "01010000001", 
		    to_sfixed(0.921514,  I, -F) when "01010000010", 
		    to_sfixed(0.920318,  I, -F) when "01010000011", 
		    to_sfixed(0.919114,  I, -F) when "01010000100", 
		    to_sfixed(0.917901,  I, -F) when "01010000101", 
		    to_sfixed(0.916679,  I, -F) when "01010000110", 
		    to_sfixed(0.915449,  I, -F) when "01010000111", 
		    to_sfixed(0.914210,  I, -F) when "01010001000", 
		    to_sfixed(0.912962,  I, -F) when "01010001001", 
		    to_sfixed(0.911706,  I, -F) when "01010001010", 
		    to_sfixed(0.910441,  I, -F) when "01010001011", 
		    to_sfixed(0.909168,  I, -F) when "01010001100", 
		    to_sfixed(0.907886,  I, -F) when "01010001101", 
		    to_sfixed(0.906596,  I, -F) when "01010001110", 
		    to_sfixed(0.905297,  I, -F) when "01010001111", 
		    to_sfixed(0.903989,  I, -F) when "01010010000", 
		    to_sfixed(0.902673,  I, -F) when "01010010001", 
		    to_sfixed(0.901349,  I, -F) when "01010010010", 
		    to_sfixed(0.900016,  I, -F) when "01010010011", 
		    to_sfixed(0.898674,  I, -F) when "01010010100", 
		    to_sfixed(0.897325,  I, -F) when "01010010101", 
		    to_sfixed(0.895966,  I, -F) when "01010010110", 
		    to_sfixed(0.894599,  I, -F) when "01010010111", 
		    to_sfixed(0.893224,  I, -F) when "01010011000", 
		    to_sfixed(0.891841,  I, -F) when "01010011001", 
		    to_sfixed(0.890449,  I, -F) when "01010011010", 
		    to_sfixed(0.889048,  I, -F) when "01010011011", 
		    to_sfixed(0.887640,  I, -F) when "01010011100", 
		    to_sfixed(0.886223,  I, -F) when "01010011101", 
		    to_sfixed(0.884797,  I, -F) when "01010011110", 
		    to_sfixed(0.883363,  I, -F) when "01010011111", 
		    to_sfixed(0.881921,  I, -F) when "01010100000", 
		    to_sfixed(0.880471,  I, -F) when "01010100001", 
		    to_sfixed(0.879012,  I, -F) when "01010100010", 
		    to_sfixed(0.877545,  I, -F) when "01010100011", 
		    to_sfixed(0.876070,  I, -F) when "01010100100", 
		    to_sfixed(0.874587,  I, -F) when "01010100101", 
		    to_sfixed(0.873095,  I, -F) when "01010100110", 
		    to_sfixed(0.871595,  I, -F) when "01010100111", 
		    to_sfixed(0.870087,  I, -F) when "01010101000", 
		    to_sfixed(0.868571,  I, -F) when "01010101001", 
		    to_sfixed(0.867046,  I, -F) when "01010101010", 
		    to_sfixed(0.865514,  I, -F) when "01010101011", 
		    to_sfixed(0.863973,  I, -F) when "01010101100", 
		    to_sfixed(0.862424,  I, -F) when "01010101101", 
		    to_sfixed(0.860867,  I, -F) when "01010101110", 
		    to_sfixed(0.859302,  I, -F) when "01010101111", 
		    to_sfixed(0.857729,  I, -F) when "01010110000", 
		    to_sfixed(0.856147,  I, -F) when "01010110001", 
		    to_sfixed(0.854558,  I, -F) when "01010110010", 
		    to_sfixed(0.852961,  I, -F) when "01010110011", 
		    to_sfixed(0.851355,  I, -F) when "01010110100", 
		    to_sfixed(0.849742,  I, -F) when "01010110101", 
		    to_sfixed(0.848120,  I, -F) when "01010110110", 
		    to_sfixed(0.846491,  I, -F) when "01010110111", 
		    to_sfixed(0.844854,  I, -F) when "01010111000", 
		    to_sfixed(0.843208,  I, -F) when "01010111001", 
		    to_sfixed(0.841555,  I, -F) when "01010111010", 
		    to_sfixed(0.839894,  I, -F) when "01010111011", 
		    to_sfixed(0.838225,  I, -F) when "01010111100", 
		    to_sfixed(0.836548,  I, -F) when "01010111101", 
		    to_sfixed(0.834863,  I, -F) when "01010111110", 
		    to_sfixed(0.833170,  I, -F) when "01010111111", 
		    to_sfixed(0.831470,  I, -F) when "01011000000", 
		    to_sfixed(0.829761,  I, -F) when "01011000001", 
		    to_sfixed(0.828045,  I, -F) when "01011000010", 
		    to_sfixed(0.826321,  I, -F) when "01011000011", 
		    to_sfixed(0.824589,  I, -F) when "01011000100", 
		    to_sfixed(0.822850,  I, -F) when "01011000101", 
		    to_sfixed(0.821103,  I, -F) when "01011000110", 
		    to_sfixed(0.819348,  I, -F) when "01011000111", 
		    to_sfixed(0.817585,  I, -F) when "01011001000", 
		    to_sfixed(0.815814,  I, -F) when "01011001001", 
		    to_sfixed(0.814036,  I, -F) when "01011001010", 
		    to_sfixed(0.812251,  I, -F) when "01011001011", 
		    to_sfixed(0.810457,  I, -F) when "01011001100", 
		    to_sfixed(0.808656,  I, -F) when "01011001101", 
		    to_sfixed(0.806848,  I, -F) when "01011001110", 
		    to_sfixed(0.805031,  I, -F) when "01011001111", 
		    to_sfixed(0.803208,  I, -F) when "01011010000", 
		    to_sfixed(0.801376,  I, -F) when "01011010001", 
		    to_sfixed(0.799537,  I, -F) when "01011010010", 
		    to_sfixed(0.797691,  I, -F) when "01011010011", 
		    to_sfixed(0.795837,  I, -F) when "01011010100", 
		    to_sfixed(0.793975,  I, -F) when "01011010101", 
		    to_sfixed(0.792107,  I, -F) when "01011010110", 
		    to_sfixed(0.790230,  I, -F) when "01011010111", 
		    to_sfixed(0.788346,  I, -F) when "01011011000", 
		    to_sfixed(0.786455,  I, -F) when "01011011001", 
		    to_sfixed(0.784557,  I, -F) when "01011011010", 
		    to_sfixed(0.782651,  I, -F) when "01011011011", 
		    to_sfixed(0.780737,  I, -F) when "01011011100", 
		    to_sfixed(0.778817,  I, -F) when "01011011101", 
		    to_sfixed(0.776888,  I, -F) when "01011011110", 
		    to_sfixed(0.774953,  I, -F) when "01011011111", 
		    to_sfixed(0.773010,  I, -F) when "01011100000", 
		    to_sfixed(0.771061,  I, -F) when "01011100001", 
		    to_sfixed(0.769103,  I, -F) when "01011100010", 
		    to_sfixed(0.767139,  I, -F) when "01011100011", 
		    to_sfixed(0.765167,  I, -F) when "01011100100", 
		    to_sfixed(0.763188,  I, -F) when "01011100101", 
		    to_sfixed(0.761202,  I, -F) when "01011100110", 
		    to_sfixed(0.759209,  I, -F) when "01011100111", 
		    to_sfixed(0.757209,  I, -F) when "01011101000", 
		    to_sfixed(0.755201,  I, -F) when "01011101001", 
		    to_sfixed(0.753187,  I, -F) when "01011101010", 
		    to_sfixed(0.751165,  I, -F) when "01011101011", 
		    to_sfixed(0.749136,  I, -F) when "01011101100", 
		    to_sfixed(0.747101,  I, -F) when "01011101101", 
		    to_sfixed(0.745058,  I, -F) when "01011101110", 
		    to_sfixed(0.743008,  I, -F) when "01011101111", 
		    to_sfixed(0.740951,  I, -F) when "01011110000", 
		    to_sfixed(0.738887,  I, -F) when "01011110001", 
		    to_sfixed(0.736817,  I, -F) when "01011110010", 
		    to_sfixed(0.734739,  I, -F) when "01011110011", 
		    to_sfixed(0.732654,  I, -F) when "01011110100", 
		    to_sfixed(0.730563,  I, -F) when "01011110101", 
		    to_sfixed(0.728464,  I, -F) when "01011110110", 
		    to_sfixed(0.726359,  I, -F) when "01011110111", 
		    to_sfixed(0.724247,  I, -F) when "01011111000", 
		    to_sfixed(0.722128,  I, -F) when "01011111001", 
		    to_sfixed(0.720003,  I, -F) when "01011111010", 
		    to_sfixed(0.717870,  I, -F) when "01011111011", 
		    to_sfixed(0.715731,  I, -F) when "01011111100", 
		    to_sfixed(0.713585,  I, -F) when "01011111101", 
		    to_sfixed(0.711432,  I, -F) when "01011111110", 
		    to_sfixed(0.709273,  I, -F) when "01011111111", 
		    to_sfixed(0.707107,  I, -F) when "01100000000", 
		    to_sfixed(0.704934,  I, -F) when "01100000001", 
		    to_sfixed(0.702755,  I, -F) when "01100000010", 
		    to_sfixed(0.700569,  I, -F) when "01100000011", 
		    to_sfixed(0.698376,  I, -F) when "01100000100", 
		    to_sfixed(0.696177,  I, -F) when "01100000101", 
		    to_sfixed(0.693971,  I, -F) when "01100000110", 
		    to_sfixed(0.691759,  I, -F) when "01100000111", 
		    to_sfixed(0.689541,  I, -F) when "01100001000", 
		    to_sfixed(0.687315,  I, -F) when "01100001001", 
		    to_sfixed(0.685084,  I, -F) when "01100001010", 
		    to_sfixed(0.682846,  I, -F) when "01100001011", 
		    to_sfixed(0.680601,  I, -F) when "01100001100", 
		    to_sfixed(0.678350,  I, -F) when "01100001101", 
		    to_sfixed(0.676093,  I, -F) when "01100001110", 
		    to_sfixed(0.673829,  I, -F) when "01100001111", 
		    to_sfixed(0.671559,  I, -F) when "01100010000", 
		    to_sfixed(0.669283,  I, -F) when "01100010001", 
		    to_sfixed(0.667000,  I, -F) when "01100010010", 
		    to_sfixed(0.664711,  I, -F) when "01100010011", 
		    to_sfixed(0.662416,  I, -F) when "01100010100", 
		    to_sfixed(0.660114,  I, -F) when "01100010101", 
		    to_sfixed(0.657807,  I, -F) when "01100010110", 
		    to_sfixed(0.655493,  I, -F) when "01100010111", 
		    to_sfixed(0.653173,  I, -F) when "01100011000", 
		    to_sfixed(0.650847,  I, -F) when "01100011001", 
		    to_sfixed(0.648514,  I, -F) when "01100011010", 
		    to_sfixed(0.646176,  I, -F) when "01100011011", 
		    to_sfixed(0.643832,  I, -F) when "01100011100", 
		    to_sfixed(0.641481,  I, -F) when "01100011101", 
		    to_sfixed(0.639124,  I, -F) when "01100011110", 
		    to_sfixed(0.636762,  I, -F) when "01100011111", 
		    to_sfixed(0.634393,  I, -F) when "01100100000", 
		    to_sfixed(0.632019,  I, -F) when "01100100001", 
		    to_sfixed(0.629638,  I, -F) when "01100100010", 
		    to_sfixed(0.627252,  I, -F) when "01100100011", 
		    to_sfixed(0.624859,  I, -F) when "01100100100", 
		    to_sfixed(0.622461,  I, -F) when "01100100101", 
		    to_sfixed(0.620057,  I, -F) when "01100100110", 
		    to_sfixed(0.617647,  I, -F) when "01100100111", 
		    to_sfixed(0.615232,  I, -F) when "01100101000", 
		    to_sfixed(0.612810,  I, -F) when "01100101001", 
		    to_sfixed(0.610383,  I, -F) when "01100101010", 
		    to_sfixed(0.607950,  I, -F) when "01100101011", 
		    to_sfixed(0.605511,  I, -F) when "01100101100", 
		    to_sfixed(0.603067,  I, -F) when "01100101101", 
		    to_sfixed(0.600616,  I, -F) when "01100101110", 
		    to_sfixed(0.598161,  I, -F) when "01100101111", 
		    to_sfixed(0.595699,  I, -F) when "01100110000", 
		    to_sfixed(0.593232,  I, -F) when "01100110001", 
		    to_sfixed(0.590760,  I, -F) when "01100110010", 
		    to_sfixed(0.588282,  I, -F) when "01100110011", 
		    to_sfixed(0.585798,  I, -F) when "01100110100", 
		    to_sfixed(0.583309,  I, -F) when "01100110101", 
		    to_sfixed(0.580814,  I, -F) when "01100110110", 
		    to_sfixed(0.578314,  I, -F) when "01100110111", 
		    to_sfixed(0.575808,  I, -F) when "01100111000", 
		    to_sfixed(0.573297,  I, -F) when "01100111001", 
		    to_sfixed(0.570781,  I, -F) when "01100111010", 
		    to_sfixed(0.568259,  I, -F) when "01100111011", 
		    to_sfixed(0.565732,  I, -F) when "01100111100", 
		    to_sfixed(0.563199,  I, -F) when "01100111101", 
		    to_sfixed(0.560662,  I, -F) when "01100111110", 
		    to_sfixed(0.558119,  I, -F) when "01100111111", 
		    to_sfixed(0.555570,  I, -F) when "01101000000", 
		    to_sfixed(0.553017,  I, -F) when "01101000001", 
		    to_sfixed(0.550458,  I, -F) when "01101000010", 
		    to_sfixed(0.547894,  I, -F) when "01101000011", 
		    to_sfixed(0.545325,  I, -F) when "01101000100", 
		    to_sfixed(0.542751,  I, -F) when "01101000101", 
		    to_sfixed(0.540171,  I, -F) when "01101000110", 
		    to_sfixed(0.537587,  I, -F) when "01101000111", 
		    to_sfixed(0.534998,  I, -F) when "01101001000", 
		    to_sfixed(0.532403,  I, -F) when "01101001001", 
		    to_sfixed(0.529804,  I, -F) when "01101001010", 
		    to_sfixed(0.527199,  I, -F) when "01101001011", 
		    to_sfixed(0.524590,  I, -F) when "01101001100", 
		    to_sfixed(0.521975,  I, -F) when "01101001101", 
		    to_sfixed(0.519356,  I, -F) when "01101001110", 
		    to_sfixed(0.516732,  I, -F) when "01101001111", 
		    to_sfixed(0.514103,  I, -F) when "01101010000", 
		    to_sfixed(0.511469,  I, -F) when "01101010001", 
		    to_sfixed(0.508830,  I, -F) when "01101010010", 
		    to_sfixed(0.506187,  I, -F) when "01101010011", 
		    to_sfixed(0.503538,  I, -F) when "01101010100", 
		    to_sfixed(0.500885,  I, -F) when "01101010101", 
		    to_sfixed(0.498228,  I, -F) when "01101010110", 
		    to_sfixed(0.495565,  I, -F) when "01101010111", 
		    to_sfixed(0.492898,  I, -F) when "01101011000", 
		    to_sfixed(0.490226,  I, -F) when "01101011001", 
		    to_sfixed(0.487550,  I, -F) when "01101011010", 
		    to_sfixed(0.484869,  I, -F) when "01101011011", 
		    to_sfixed(0.482184,  I, -F) when "01101011100", 
		    to_sfixed(0.479494,  I, -F) when "01101011101", 
		    to_sfixed(0.476799,  I, -F) when "01101011110", 
		    to_sfixed(0.474100,  I, -F) when "01101011111", 
		    to_sfixed(0.471397,  I, -F) when "01101100000", 
		    to_sfixed(0.468689,  I, -F) when "01101100001", 
		    to_sfixed(0.465976,  I, -F) when "01101100010", 
		    to_sfixed(0.463260,  I, -F) when "01101100011", 
		    to_sfixed(0.460539,  I, -F) when "01101100100", 
		    to_sfixed(0.457813,  I, -F) when "01101100101", 
		    to_sfixed(0.455084,  I, -F) when "01101100110", 
		    to_sfixed(0.452350,  I, -F) when "01101100111", 
		    to_sfixed(0.449611,  I, -F) when "01101101000", 
		    to_sfixed(0.446869,  I, -F) when "01101101001", 
		    to_sfixed(0.444122,  I, -F) when "01101101010", 
		    to_sfixed(0.441371,  I, -F) when "01101101011", 
		    to_sfixed(0.438616,  I, -F) when "01101101100", 
		    to_sfixed(0.435857,  I, -F) when "01101101101", 
		    to_sfixed(0.433094,  I, -F) when "01101101110", 
		    to_sfixed(0.430326,  I, -F) when "01101101111", 
		    to_sfixed(0.427555,  I, -F) when "01101110000", 
		    to_sfixed(0.424780,  I, -F) when "01101110001", 
		    to_sfixed(0.422000,  I, -F) when "01101110010", 
		    to_sfixed(0.419217,  I, -F) when "01101110011", 
		    to_sfixed(0.416430,  I, -F) when "01101110100", 
		    to_sfixed(0.413638,  I, -F) when "01101110101", 
		    to_sfixed(0.410843,  I, -F) when "01101110110", 
		    to_sfixed(0.408044,  I, -F) when "01101110111", 
		    to_sfixed(0.405241,  I, -F) when "01101111000", 
		    to_sfixed(0.402435,  I, -F) when "01101111001", 
		    to_sfixed(0.399624,  I, -F) when "01101111010", 
		    to_sfixed(0.396810,  I, -F) when "01101111011", 
		    to_sfixed(0.393992,  I, -F) when "01101111100", 
		    to_sfixed(0.391170,  I, -F) when "01101111101", 
		    to_sfixed(0.388345,  I, -F) when "01101111110", 
		    to_sfixed(0.385516,  I, -F) when "01101111111", 
		    to_sfixed(0.382683,  I, -F) when "01110000000", 
		    to_sfixed(0.379847,  I, -F) when "01110000001", 
		    to_sfixed(0.377007,  I, -F) when "01110000010", 
		    to_sfixed(0.374164,  I, -F) when "01110000011", 
		    to_sfixed(0.371317,  I, -F) when "01110000100", 
		    to_sfixed(0.368467,  I, -F) when "01110000101", 
		    to_sfixed(0.365613,  I, -F) when "01110000110", 
		    to_sfixed(0.362756,  I, -F) when "01110000111", 
		    to_sfixed(0.359895,  I, -F) when "01110001000", 
		    to_sfixed(0.357031,  I, -F) when "01110001001", 
		    to_sfixed(0.354164,  I, -F) when "01110001010", 
		    to_sfixed(0.351293,  I, -F) when "01110001011", 
		    to_sfixed(0.348419,  I, -F) when "01110001100", 
		    to_sfixed(0.345541,  I, -F) when "01110001101", 
		    to_sfixed(0.342661,  I, -F) when "01110001110", 
		    to_sfixed(0.339777,  I, -F) when "01110001111", 
		    to_sfixed(0.336890,  I, -F) when "01110010000", 
		    to_sfixed(0.334000,  I, -F) when "01110010001", 
		    to_sfixed(0.331106,  I, -F) when "01110010010", 
		    to_sfixed(0.328210,  I, -F) when "01110010011", 
		    to_sfixed(0.325310,  I, -F) when "01110010100", 
		    to_sfixed(0.322408,  I, -F) when "01110010101", 
		    to_sfixed(0.319502,  I, -F) when "01110010110", 
		    to_sfixed(0.316593,  I, -F) when "01110010111", 
		    to_sfixed(0.313682,  I, -F) when "01110011000", 
		    to_sfixed(0.310767,  I, -F) when "01110011001", 
		    to_sfixed(0.307850,  I, -F) when "01110011010", 
		    to_sfixed(0.304929,  I, -F) when "01110011011", 
		    to_sfixed(0.302006,  I, -F) when "01110011100", 
		    to_sfixed(0.299080,  I, -F) when "01110011101", 
		    to_sfixed(0.296151,  I, -F) when "01110011110", 
		    to_sfixed(0.293219,  I, -F) when "01110011111", 
		    to_sfixed(0.290285,  I, -F) when "01110100000", 
		    to_sfixed(0.287347,  I, -F) when "01110100001", 
		    to_sfixed(0.284408,  I, -F) when "01110100010", 
		    to_sfixed(0.281465,  I, -F) when "01110100011", 
		    to_sfixed(0.278520,  I, -F) when "01110100100", 
		    to_sfixed(0.275572,  I, -F) when "01110100101", 
		    to_sfixed(0.272621,  I, -F) when "01110100110", 
		    to_sfixed(0.269668,  I, -F) when "01110100111", 
		    to_sfixed(0.266713,  I, -F) when "01110101000", 
		    to_sfixed(0.263755,  I, -F) when "01110101001", 
		    to_sfixed(0.260794,  I, -F) when "01110101010", 
		    to_sfixed(0.257831,  I, -F) when "01110101011", 
		    to_sfixed(0.254866,  I, -F) when "01110101100", 
		    to_sfixed(0.251898,  I, -F) when "01110101101", 
		    to_sfixed(0.248928,  I, -F) when "01110101110", 
		    to_sfixed(0.245955,  I, -F) when "01110101111", 
		    to_sfixed(0.242980,  I, -F) when "01110110000", 
		    to_sfixed(0.240003,  I, -F) when "01110110001", 
		    to_sfixed(0.237024,  I, -F) when "01110110010", 
		    to_sfixed(0.234042,  I, -F) when "01110110011", 
		    to_sfixed(0.231058,  I, -F) when "01110110100", 
		    to_sfixed(0.228072,  I, -F) when "01110110101", 
		    to_sfixed(0.225084,  I, -F) when "01110110110", 
		    to_sfixed(0.222094,  I, -F) when "01110110111", 
		    to_sfixed(0.219101,  I, -F) when "01110111000", 
		    to_sfixed(0.216107,  I, -F) when "01110111001", 
		    to_sfixed(0.213110,  I, -F) when "01110111010", 
		    to_sfixed(0.210112,  I, -F) when "01110111011", 
		    to_sfixed(0.207111,  I, -F) when "01110111100", 
		    to_sfixed(0.204109,  I, -F) when "01110111101", 
		    to_sfixed(0.201105,  I, -F) when "01110111110", 
		    to_sfixed(0.198098,  I, -F) when "01110111111", 
		    to_sfixed(0.195090,  I, -F) when "01111000000", 
		    to_sfixed(0.192080,  I, -F) when "01111000001", 
		    to_sfixed(0.189069,  I, -F) when "01111000010", 
		    to_sfixed(0.186055,  I, -F) when "01111000011", 
		    to_sfixed(0.183040,  I, -F) when "01111000100", 
		    to_sfixed(0.180023,  I, -F) when "01111000101", 
		    to_sfixed(0.177004,  I, -F) when "01111000110", 
		    to_sfixed(0.173984,  I, -F) when "01111000111", 
		    to_sfixed(0.170962,  I, -F) when "01111001000", 
		    to_sfixed(0.167938,  I, -F) when "01111001001", 
		    to_sfixed(0.164913,  I, -F) when "01111001010", 
		    to_sfixed(0.161886,  I, -F) when "01111001011", 
		    to_sfixed(0.158858,  I, -F) when "01111001100", 
		    to_sfixed(0.155828,  I, -F) when "01111001101", 
		    to_sfixed(0.152797,  I, -F) when "01111001110", 
		    to_sfixed(0.149765,  I, -F) when "01111001111", 
		    to_sfixed(0.146730,  I, -F) when "01111010000", 
		    to_sfixed(0.143695,  I, -F) when "01111010001", 
		    to_sfixed(0.140658,  I, -F) when "01111010010", 
		    to_sfixed(0.137620,  I, -F) when "01111010011", 
		    to_sfixed(0.134581,  I, -F) when "01111010100", 
		    to_sfixed(0.131540,  I, -F) when "01111010101", 
		    to_sfixed(0.128498,  I, -F) when "01111010110", 
		    to_sfixed(0.125455,  I, -F) when "01111010111", 
		    to_sfixed(0.122411,  I, -F) when "01111011000", 
		    to_sfixed(0.119365,  I, -F) when "01111011001", 
		    to_sfixed(0.116319,  I, -F) when "01111011010", 
		    to_sfixed(0.113271,  I, -F) when "01111011011", 
		    to_sfixed(0.110222,  I, -F) when "01111011100", 
		    to_sfixed(0.107172,  I, -F) when "01111011101", 
		    to_sfixed(0.104122,  I, -F) when "01111011110", 
		    to_sfixed(0.101070,  I, -F) when "01111011111", 
		    to_sfixed(0.098017,  I, -F) when "01111100000", 
		    to_sfixed(0.094963,  I, -F) when "01111100001", 
		    to_sfixed(0.091909,  I, -F) when "01111100010", 
		    to_sfixed(0.088854,  I, -F) when "01111100011", 
		    to_sfixed(0.085797,  I, -F) when "01111100100", 
		    to_sfixed(0.082740,  I, -F) when "01111100101", 
		    to_sfixed(0.079682,  I, -F) when "01111100110", 
		    to_sfixed(0.076624,  I, -F) when "01111100111", 
		    to_sfixed(0.073565,  I, -F) when "01111101000", 
		    to_sfixed(0.070505,  I, -F) when "01111101001", 
		    to_sfixed(0.067444,  I, -F) when "01111101010", 
		    to_sfixed(0.064383,  I, -F) when "01111101011", 
		    to_sfixed(0.061321,  I, -F) when "01111101100", 
		    to_sfixed(0.058258,  I, -F) when "01111101101", 
		    to_sfixed(0.055195,  I, -F) when "01111101110", 
		    to_sfixed(0.052132,  I, -F) when "01111101111", 
		    to_sfixed(0.049068,  I, -F) when "01111110000", 
		    to_sfixed(0.046003,  I, -F) when "01111110001", 
		    to_sfixed(0.042938,  I, -F) when "01111110010", 
		    to_sfixed(0.039873,  I, -F) when "01111110011", 
		    to_sfixed(0.036807,  I, -F) when "01111110100", 
		    to_sfixed(0.033741,  I, -F) when "01111110101", 
		    to_sfixed(0.030675,  I, -F) when "01111110110", 
		    to_sfixed(0.027608,  I, -F) when "01111110111", 
		    to_sfixed(0.024541,  I, -F) when "01111111000", 
		    to_sfixed(0.021474,  I, -F) when "01111111001", 
		    to_sfixed(0.018407,  I, -F) when "01111111010", 
		    to_sfixed(0.015339,  I, -F) when "01111111011", 
		    to_sfixed(0.012272,  I, -F) when "01111111100", 
		    to_sfixed(0.009204,  I, -F) when "01111111101", 
		    to_sfixed(0.006136,  I, -F) when "01111111110", 
		    to_sfixed(0.003068,  I, -F) when "01111111111", 
		    to_sfixed(0.000000,  I, -F) when "10000000000", 
		    to_sfixed(-0.003068,  I, -F) when "10000000001", 
		    to_sfixed(-0.006136,  I, -F) when "10000000010", 
		    to_sfixed(-0.009204,  I, -F) when "10000000011", 
		    to_sfixed(-0.012272,  I, -F) when "10000000100", 
		    to_sfixed(-0.015339,  I, -F) when "10000000101", 
		    to_sfixed(-0.018407,  I, -F) when "10000000110", 
		    to_sfixed(-0.021474,  I, -F) when "10000000111", 
		    to_sfixed(-0.024541,  I, -F) when "10000001000", 
		    to_sfixed(-0.027608,  I, -F) when "10000001001", 
		    to_sfixed(-0.030675,  I, -F) when "10000001010", 
		    to_sfixed(-0.033741,  I, -F) when "10000001011", 
		    to_sfixed(-0.036807,  I, -F) when "10000001100", 
		    to_sfixed(-0.039873,  I, -F) when "10000001101", 
		    to_sfixed(-0.042938,  I, -F) when "10000001110", 
		    to_sfixed(-0.046003,  I, -F) when "10000001111", 
		    to_sfixed(-0.049068,  I, -F) when "10000010000", 
		    to_sfixed(-0.052132,  I, -F) when "10000010001", 
		    to_sfixed(-0.055195,  I, -F) when "10000010010", 
		    to_sfixed(-0.058258,  I, -F) when "10000010011", 
		    to_sfixed(-0.061321,  I, -F) when "10000010100", 
		    to_sfixed(-0.064383,  I, -F) when "10000010101", 
		    to_sfixed(-0.067444,  I, -F) when "10000010110", 
		    to_sfixed(-0.070505,  I, -F) when "10000010111", 
		    to_sfixed(-0.073565,  I, -F) when "10000011000", 
		    to_sfixed(-0.076624,  I, -F) when "10000011001", 
		    to_sfixed(-0.079682,  I, -F) when "10000011010", 
		    to_sfixed(-0.082740,  I, -F) when "10000011011", 
		    to_sfixed(-0.085797,  I, -F) when "10000011100", 
		    to_sfixed(-0.088854,  I, -F) when "10000011101", 
		    to_sfixed(-0.091909,  I, -F) when "10000011110", 
		    to_sfixed(-0.094963,  I, -F) when "10000011111", 
		    to_sfixed(-0.098017,  I, -F) when "10000100000", 
		    to_sfixed(-0.101070,  I, -F) when "10000100001", 
		    to_sfixed(-0.104122,  I, -F) when "10000100010", 
		    to_sfixed(-0.107172,  I, -F) when "10000100011", 
		    to_sfixed(-0.110222,  I, -F) when "10000100100", 
		    to_sfixed(-0.113271,  I, -F) when "10000100101", 
		    to_sfixed(-0.116319,  I, -F) when "10000100110", 
		    to_sfixed(-0.119365,  I, -F) when "10000100111", 
		    to_sfixed(-0.122411,  I, -F) when "10000101000", 
		    to_sfixed(-0.125455,  I, -F) when "10000101001", 
		    to_sfixed(-0.128498,  I, -F) when "10000101010", 
		    to_sfixed(-0.131540,  I, -F) when "10000101011", 
		    to_sfixed(-0.134581,  I, -F) when "10000101100", 
		    to_sfixed(-0.137620,  I, -F) when "10000101101", 
		    to_sfixed(-0.140658,  I, -F) when "10000101110", 
		    to_sfixed(-0.143695,  I, -F) when "10000101111", 
		    to_sfixed(-0.146730,  I, -F) when "10000110000", 
		    to_sfixed(-0.149765,  I, -F) when "10000110001", 
		    to_sfixed(-0.152797,  I, -F) when "10000110010", 
		    to_sfixed(-0.155828,  I, -F) when "10000110011", 
		    to_sfixed(-0.158858,  I, -F) when "10000110100", 
		    to_sfixed(-0.161886,  I, -F) when "10000110101", 
		    to_sfixed(-0.164913,  I, -F) when "10000110110", 
		    to_sfixed(-0.167938,  I, -F) when "10000110111", 
		    to_sfixed(-0.170962,  I, -F) when "10000111000", 
		    to_sfixed(-0.173984,  I, -F) when "10000111001", 
		    to_sfixed(-0.177004,  I, -F) when "10000111010", 
		    to_sfixed(-0.180023,  I, -F) when "10000111011", 
		    to_sfixed(-0.183040,  I, -F) when "10000111100", 
		    to_sfixed(-0.186055,  I, -F) when "10000111101", 
		    to_sfixed(-0.189069,  I, -F) when "10000111110", 
		    to_sfixed(-0.192080,  I, -F) when "10000111111", 
		    to_sfixed(-0.195090,  I, -F) when "10001000000", 
		    to_sfixed(-0.198098,  I, -F) when "10001000001", 
		    to_sfixed(-0.201105,  I, -F) when "10001000010", 
		    to_sfixed(-0.204109,  I, -F) when "10001000011", 
		    to_sfixed(-0.207111,  I, -F) when "10001000100", 
		    to_sfixed(-0.210112,  I, -F) when "10001000101", 
		    to_sfixed(-0.213110,  I, -F) when "10001000110", 
		    to_sfixed(-0.216107,  I, -F) when "10001000111", 
		    to_sfixed(-0.219101,  I, -F) when "10001001000", 
		    to_sfixed(-0.222094,  I, -F) when "10001001001", 
		    to_sfixed(-0.225084,  I, -F) when "10001001010", 
		    to_sfixed(-0.228072,  I, -F) when "10001001011", 
		    to_sfixed(-0.231058,  I, -F) when "10001001100", 
		    to_sfixed(-0.234042,  I, -F) when "10001001101", 
		    to_sfixed(-0.237024,  I, -F) when "10001001110", 
		    to_sfixed(-0.240003,  I, -F) when "10001001111", 
		    to_sfixed(-0.242980,  I, -F) when "10001010000", 
		    to_sfixed(-0.245955,  I, -F) when "10001010001", 
		    to_sfixed(-0.248928,  I, -F) when "10001010010", 
		    to_sfixed(-0.251898,  I, -F) when "10001010011", 
		    to_sfixed(-0.254866,  I, -F) when "10001010100", 
		    to_sfixed(-0.257831,  I, -F) when "10001010101", 
		    to_sfixed(-0.260794,  I, -F) when "10001010110", 
		    to_sfixed(-0.263755,  I, -F) when "10001010111", 
		    to_sfixed(-0.266713,  I, -F) when "10001011000", 
		    to_sfixed(-0.269668,  I, -F) when "10001011001", 
		    to_sfixed(-0.272621,  I, -F) when "10001011010", 
		    to_sfixed(-0.275572,  I, -F) when "10001011011", 
		    to_sfixed(-0.278520,  I, -F) when "10001011100", 
		    to_sfixed(-0.281465,  I, -F) when "10001011101", 
		    to_sfixed(-0.284408,  I, -F) when "10001011110", 
		    to_sfixed(-0.287347,  I, -F) when "10001011111", 
		    to_sfixed(-0.290285,  I, -F) when "10001100000", 
		    to_sfixed(-0.293219,  I, -F) when "10001100001", 
		    to_sfixed(-0.296151,  I, -F) when "10001100010", 
		    to_sfixed(-0.299080,  I, -F) when "10001100011", 
		    to_sfixed(-0.302006,  I, -F) when "10001100100", 
		    to_sfixed(-0.304929,  I, -F) when "10001100101", 
		    to_sfixed(-0.307850,  I, -F) when "10001100110", 
		    to_sfixed(-0.310767,  I, -F) when "10001100111", 
		    to_sfixed(-0.313682,  I, -F) when "10001101000", 
		    to_sfixed(-0.316593,  I, -F) when "10001101001", 
		    to_sfixed(-0.319502,  I, -F) when "10001101010", 
		    to_sfixed(-0.322408,  I, -F) when "10001101011", 
		    to_sfixed(-0.325310,  I, -F) when "10001101100", 
		    to_sfixed(-0.328210,  I, -F) when "10001101101", 
		    to_sfixed(-0.331106,  I, -F) when "10001101110", 
		    to_sfixed(-0.334000,  I, -F) when "10001101111", 
		    to_sfixed(-0.336890,  I, -F) when "10001110000", 
		    to_sfixed(-0.339777,  I, -F) when "10001110001", 
		    to_sfixed(-0.342661,  I, -F) when "10001110010", 
		    to_sfixed(-0.345541,  I, -F) when "10001110011", 
		    to_sfixed(-0.348419,  I, -F) when "10001110100", 
		    to_sfixed(-0.351293,  I, -F) when "10001110101", 
		    to_sfixed(-0.354164,  I, -F) when "10001110110", 
		    to_sfixed(-0.357031,  I, -F) when "10001110111", 
		    to_sfixed(-0.359895,  I, -F) when "10001111000", 
		    to_sfixed(-0.362756,  I, -F) when "10001111001", 
		    to_sfixed(-0.365613,  I, -F) when "10001111010", 
		    to_sfixed(-0.368467,  I, -F) when "10001111011", 
		    to_sfixed(-0.371317,  I, -F) when "10001111100", 
		    to_sfixed(-0.374164,  I, -F) when "10001111101", 
		    to_sfixed(-0.377007,  I, -F) when "10001111110", 
		    to_sfixed(-0.379847,  I, -F) when "10001111111", 
		    to_sfixed(-0.382683,  I, -F) when "10010000000", 
		    to_sfixed(-0.385516,  I, -F) when "10010000001", 
		    to_sfixed(-0.388345,  I, -F) when "10010000010", 
		    to_sfixed(-0.391170,  I, -F) when "10010000011", 
		    to_sfixed(-0.393992,  I, -F) when "10010000100", 
		    to_sfixed(-0.396810,  I, -F) when "10010000101", 
		    to_sfixed(-0.399624,  I, -F) when "10010000110", 
		    to_sfixed(-0.402435,  I, -F) when "10010000111", 
		    to_sfixed(-0.405241,  I, -F) when "10010001000", 
		    to_sfixed(-0.408044,  I, -F) when "10010001001", 
		    to_sfixed(-0.410843,  I, -F) when "10010001010", 
		    to_sfixed(-0.413638,  I, -F) when "10010001011", 
		    to_sfixed(-0.416430,  I, -F) when "10010001100", 
		    to_sfixed(-0.419217,  I, -F) when "10010001101", 
		    to_sfixed(-0.422000,  I, -F) when "10010001110", 
		    to_sfixed(-0.424780,  I, -F) when "10010001111", 
		    to_sfixed(-0.427555,  I, -F) when "10010010000", 
		    to_sfixed(-0.430326,  I, -F) when "10010010001", 
		    to_sfixed(-0.433094,  I, -F) when "10010010010", 
		    to_sfixed(-0.435857,  I, -F) when "10010010011", 
		    to_sfixed(-0.438616,  I, -F) when "10010010100", 
		    to_sfixed(-0.441371,  I, -F) when "10010010101", 
		    to_sfixed(-0.444122,  I, -F) when "10010010110", 
		    to_sfixed(-0.446869,  I, -F) when "10010010111", 
		    to_sfixed(-0.449611,  I, -F) when "10010011000", 
		    to_sfixed(-0.452350,  I, -F) when "10010011001", 
		    to_sfixed(-0.455084,  I, -F) when "10010011010", 
		    to_sfixed(-0.457813,  I, -F) when "10010011011", 
		    to_sfixed(-0.460539,  I, -F) when "10010011100", 
		    to_sfixed(-0.463260,  I, -F) when "10010011101", 
		    to_sfixed(-0.465976,  I, -F) when "10010011110", 
		    to_sfixed(-0.468689,  I, -F) when "10010011111", 
		    to_sfixed(-0.471397,  I, -F) when "10010100000", 
		    to_sfixed(-0.474100,  I, -F) when "10010100001", 
		    to_sfixed(-0.476799,  I, -F) when "10010100010", 
		    to_sfixed(-0.479494,  I, -F) when "10010100011", 
		    to_sfixed(-0.482184,  I, -F) when "10010100100", 
		    to_sfixed(-0.484869,  I, -F) when "10010100101", 
		    to_sfixed(-0.487550,  I, -F) when "10010100110", 
		    to_sfixed(-0.490226,  I, -F) when "10010100111", 
		    to_sfixed(-0.492898,  I, -F) when "10010101000", 
		    to_sfixed(-0.495565,  I, -F) when "10010101001", 
		    to_sfixed(-0.498228,  I, -F) when "10010101010", 
		    to_sfixed(-0.500885,  I, -F) when "10010101011", 
		    to_sfixed(-0.503538,  I, -F) when "10010101100", 
		    to_sfixed(-0.506187,  I, -F) when "10010101101", 
		    to_sfixed(-0.508830,  I, -F) when "10010101110", 
		    to_sfixed(-0.511469,  I, -F) when "10010101111", 
		    to_sfixed(-0.514103,  I, -F) when "10010110000", 
		    to_sfixed(-0.516732,  I, -F) when "10010110001", 
		    to_sfixed(-0.519356,  I, -F) when "10010110010", 
		    to_sfixed(-0.521975,  I, -F) when "10010110011", 
		    to_sfixed(-0.524590,  I, -F) when "10010110100", 
		    to_sfixed(-0.527199,  I, -F) when "10010110101", 
		    to_sfixed(-0.529804,  I, -F) when "10010110110", 
		    to_sfixed(-0.532403,  I, -F) when "10010110111", 
		    to_sfixed(-0.534998,  I, -F) when "10010111000", 
		    to_sfixed(-0.537587,  I, -F) when "10010111001", 
		    to_sfixed(-0.540171,  I, -F) when "10010111010", 
		    to_sfixed(-0.542751,  I, -F) when "10010111011", 
		    to_sfixed(-0.545325,  I, -F) when "10010111100", 
		    to_sfixed(-0.547894,  I, -F) when "10010111101", 
		    to_sfixed(-0.550458,  I, -F) when "10010111110", 
		    to_sfixed(-0.553017,  I, -F) when "10010111111", 
		    to_sfixed(-0.555570,  I, -F) when "10011000000", 
		    to_sfixed(-0.558119,  I, -F) when "10011000001", 
		    to_sfixed(-0.560662,  I, -F) when "10011000010", 
		    to_sfixed(-0.563199,  I, -F) when "10011000011", 
		    to_sfixed(-0.565732,  I, -F) when "10011000100", 
		    to_sfixed(-0.568259,  I, -F) when "10011000101", 
		    to_sfixed(-0.570781,  I, -F) when "10011000110", 
		    to_sfixed(-0.573297,  I, -F) when "10011000111", 
		    to_sfixed(-0.575808,  I, -F) when "10011001000", 
		    to_sfixed(-0.578314,  I, -F) when "10011001001", 
		    to_sfixed(-0.580814,  I, -F) when "10011001010", 
		    to_sfixed(-0.583309,  I, -F) when "10011001011", 
		    to_sfixed(-0.585798,  I, -F) when "10011001100", 
		    to_sfixed(-0.588282,  I, -F) when "10011001101", 
		    to_sfixed(-0.590760,  I, -F) when "10011001110", 
		    to_sfixed(-0.593232,  I, -F) when "10011001111", 
		    to_sfixed(-0.595699,  I, -F) when "10011010000", 
		    to_sfixed(-0.598161,  I, -F) when "10011010001", 
		    to_sfixed(-0.600616,  I, -F) when "10011010010", 
		    to_sfixed(-0.603067,  I, -F) when "10011010011", 
		    to_sfixed(-0.605511,  I, -F) when "10011010100", 
		    to_sfixed(-0.607950,  I, -F) when "10011010101", 
		    to_sfixed(-0.610383,  I, -F) when "10011010110", 
		    to_sfixed(-0.612810,  I, -F) when "10011010111", 
		    to_sfixed(-0.615232,  I, -F) when "10011011000", 
		    to_sfixed(-0.617647,  I, -F) when "10011011001", 
		    to_sfixed(-0.620057,  I, -F) when "10011011010", 
		    to_sfixed(-0.622461,  I, -F) when "10011011011", 
		    to_sfixed(-0.624859,  I, -F) when "10011011100", 
		    to_sfixed(-0.627252,  I, -F) when "10011011101", 
		    to_sfixed(-0.629638,  I, -F) when "10011011110", 
		    to_sfixed(-0.632019,  I, -F) when "10011011111", 
		    to_sfixed(-0.634393,  I, -F) when "10011100000", 
		    to_sfixed(-0.636762,  I, -F) when "10011100001", 
		    to_sfixed(-0.639124,  I, -F) when "10011100010", 
		    to_sfixed(-0.641481,  I, -F) when "10011100011", 
		    to_sfixed(-0.643832,  I, -F) when "10011100100", 
		    to_sfixed(-0.646176,  I, -F) when "10011100101", 
		    to_sfixed(-0.648514,  I, -F) when "10011100110", 
		    to_sfixed(-0.650847,  I, -F) when "10011100111", 
		    to_sfixed(-0.653173,  I, -F) when "10011101000", 
		    to_sfixed(-0.655493,  I, -F) when "10011101001", 
		    to_sfixed(-0.657807,  I, -F) when "10011101010", 
		    to_sfixed(-0.660114,  I, -F) when "10011101011", 
		    to_sfixed(-0.662416,  I, -F) when "10011101100", 
		    to_sfixed(-0.664711,  I, -F) when "10011101101", 
		    to_sfixed(-0.667000,  I, -F) when "10011101110", 
		    to_sfixed(-0.669283,  I, -F) when "10011101111", 
		    to_sfixed(-0.671559,  I, -F) when "10011110000", 
		    to_sfixed(-0.673829,  I, -F) when "10011110001", 
		    to_sfixed(-0.676093,  I, -F) when "10011110010", 
		    to_sfixed(-0.678350,  I, -F) when "10011110011", 
		    to_sfixed(-0.680601,  I, -F) when "10011110100", 
		    to_sfixed(-0.682846,  I, -F) when "10011110101", 
		    to_sfixed(-0.685084,  I, -F) when "10011110110", 
		    to_sfixed(-0.687315,  I, -F) when "10011110111", 
		    to_sfixed(-0.689541,  I, -F) when "10011111000", 
		    to_sfixed(-0.691759,  I, -F) when "10011111001", 
		    to_sfixed(-0.693971,  I, -F) when "10011111010", 
		    to_sfixed(-0.696177,  I, -F) when "10011111011", 
		    to_sfixed(-0.698376,  I, -F) when "10011111100", 
		    to_sfixed(-0.700569,  I, -F) when "10011111101", 
		    to_sfixed(-0.702755,  I, -F) when "10011111110", 
		    to_sfixed(-0.704934,  I, -F) when "10011111111", 
		    to_sfixed(-0.707107,  I, -F) when "10100000000", 
		    to_sfixed(-0.709273,  I, -F) when "10100000001", 
		    to_sfixed(-0.711432,  I, -F) when "10100000010", 
		    to_sfixed(-0.713585,  I, -F) when "10100000011", 
		    to_sfixed(-0.715731,  I, -F) when "10100000100", 
		    to_sfixed(-0.717870,  I, -F) when "10100000101", 
		    to_sfixed(-0.720003,  I, -F) when "10100000110", 
		    to_sfixed(-0.722128,  I, -F) when "10100000111", 
		    to_sfixed(-0.724247,  I, -F) when "10100001000", 
		    to_sfixed(-0.726359,  I, -F) when "10100001001", 
		    to_sfixed(-0.728464,  I, -F) when "10100001010", 
		    to_sfixed(-0.730563,  I, -F) when "10100001011", 
		    to_sfixed(-0.732654,  I, -F) when "10100001100", 
		    to_sfixed(-0.734739,  I, -F) when "10100001101", 
		    to_sfixed(-0.736817,  I, -F) when "10100001110", 
		    to_sfixed(-0.738887,  I, -F) when "10100001111", 
		    to_sfixed(-0.740951,  I, -F) when "10100010000", 
		    to_sfixed(-0.743008,  I, -F) when "10100010001", 
		    to_sfixed(-0.745058,  I, -F) when "10100010010", 
		    to_sfixed(-0.747101,  I, -F) when "10100010011", 
		    to_sfixed(-0.749136,  I, -F) when "10100010100", 
		    to_sfixed(-0.751165,  I, -F) when "10100010101", 
		    to_sfixed(-0.753187,  I, -F) when "10100010110", 
		    to_sfixed(-0.755201,  I, -F) when "10100010111", 
		    to_sfixed(-0.757209,  I, -F) when "10100011000", 
		    to_sfixed(-0.759209,  I, -F) when "10100011001", 
		    to_sfixed(-0.761202,  I, -F) when "10100011010", 
		    to_sfixed(-0.763188,  I, -F) when "10100011011", 
		    to_sfixed(-0.765167,  I, -F) when "10100011100", 
		    to_sfixed(-0.767139,  I, -F) when "10100011101", 
		    to_sfixed(-0.769103,  I, -F) when "10100011110", 
		    to_sfixed(-0.771061,  I, -F) when "10100011111", 
		    to_sfixed(-0.773010,  I, -F) when "10100100000", 
		    to_sfixed(-0.774953,  I, -F) when "10100100001", 
		    to_sfixed(-0.776888,  I, -F) when "10100100010", 
		    to_sfixed(-0.778817,  I, -F) when "10100100011", 
		    to_sfixed(-0.780737,  I, -F) when "10100100100", 
		    to_sfixed(-0.782651,  I, -F) when "10100100101", 
		    to_sfixed(-0.784557,  I, -F) when "10100100110", 
		    to_sfixed(-0.786455,  I, -F) when "10100100111", 
		    to_sfixed(-0.788346,  I, -F) when "10100101000", 
		    to_sfixed(-0.790230,  I, -F) when "10100101001", 
		    to_sfixed(-0.792107,  I, -F) when "10100101010", 
		    to_sfixed(-0.793975,  I, -F) when "10100101011", 
		    to_sfixed(-0.795837,  I, -F) when "10100101100", 
		    to_sfixed(-0.797691,  I, -F) when "10100101101", 
		    to_sfixed(-0.799537,  I, -F) when "10100101110", 
		    to_sfixed(-0.801376,  I, -F) when "10100101111", 
		    to_sfixed(-0.803208,  I, -F) when "10100110000", 
		    to_sfixed(-0.805031,  I, -F) when "10100110001", 
		    to_sfixed(-0.806848,  I, -F) when "10100110010", 
		    to_sfixed(-0.808656,  I, -F) when "10100110011", 
		    to_sfixed(-0.810457,  I, -F) when "10100110100", 
		    to_sfixed(-0.812251,  I, -F) when "10100110101", 
		    to_sfixed(-0.814036,  I, -F) when "10100110110", 
		    to_sfixed(-0.815814,  I, -F) when "10100110111", 
		    to_sfixed(-0.817585,  I, -F) when "10100111000", 
		    to_sfixed(-0.819348,  I, -F) when "10100111001", 
		    to_sfixed(-0.821103,  I, -F) when "10100111010", 
		    to_sfixed(-0.822850,  I, -F) when "10100111011", 
		    to_sfixed(-0.824589,  I, -F) when "10100111100", 
		    to_sfixed(-0.826321,  I, -F) when "10100111101", 
		    to_sfixed(-0.828045,  I, -F) when "10100111110", 
		    to_sfixed(-0.829761,  I, -F) when "10100111111", 
		    to_sfixed(-0.831470,  I, -F) when "10101000000", 
		    to_sfixed(-0.833170,  I, -F) when "10101000001", 
		    to_sfixed(-0.834863,  I, -F) when "10101000010", 
		    to_sfixed(-0.836548,  I, -F) when "10101000011", 
		    to_sfixed(-0.838225,  I, -F) when "10101000100", 
		    to_sfixed(-0.839894,  I, -F) when "10101000101", 
		    to_sfixed(-0.841555,  I, -F) when "10101000110", 
		    to_sfixed(-0.843208,  I, -F) when "10101000111", 
		    to_sfixed(-0.844854,  I, -F) when "10101001000", 
		    to_sfixed(-0.846491,  I, -F) when "10101001001", 
		    to_sfixed(-0.848120,  I, -F) when "10101001010", 
		    to_sfixed(-0.849742,  I, -F) when "10101001011", 
		    to_sfixed(-0.851355,  I, -F) when "10101001100", 
		    to_sfixed(-0.852961,  I, -F) when "10101001101", 
		    to_sfixed(-0.854558,  I, -F) when "10101001110", 
		    to_sfixed(-0.856147,  I, -F) when "10101001111", 
		    to_sfixed(-0.857729,  I, -F) when "10101010000", 
		    to_sfixed(-0.859302,  I, -F) when "10101010001", 
		    to_sfixed(-0.860867,  I, -F) when "10101010010", 
		    to_sfixed(-0.862424,  I, -F) when "10101010011", 
		    to_sfixed(-0.863973,  I, -F) when "10101010100", 
		    to_sfixed(-0.865514,  I, -F) when "10101010101", 
		    to_sfixed(-0.867046,  I, -F) when "10101010110", 
		    to_sfixed(-0.868571,  I, -F) when "10101010111", 
		    to_sfixed(-0.870087,  I, -F) when "10101011000", 
		    to_sfixed(-0.871595,  I, -F) when "10101011001", 
		    to_sfixed(-0.873095,  I, -F) when "10101011010", 
		    to_sfixed(-0.874587,  I, -F) when "10101011011", 
		    to_sfixed(-0.876070,  I, -F) when "10101011100", 
		    to_sfixed(-0.877545,  I, -F) when "10101011101", 
		    to_sfixed(-0.879012,  I, -F) when "10101011110", 
		    to_sfixed(-0.880471,  I, -F) when "10101011111", 
		    to_sfixed(-0.881921,  I, -F) when "10101100000", 
		    to_sfixed(-0.883363,  I, -F) when "10101100001", 
		    to_sfixed(-0.884797,  I, -F) when "10101100010", 
		    to_sfixed(-0.886223,  I, -F) when "10101100011", 
		    to_sfixed(-0.887640,  I, -F) when "10101100100", 
		    to_sfixed(-0.889048,  I, -F) when "10101100101", 
		    to_sfixed(-0.890449,  I, -F) when "10101100110", 
		    to_sfixed(-0.891841,  I, -F) when "10101100111", 
		    to_sfixed(-0.893224,  I, -F) when "10101101000", 
		    to_sfixed(-0.894599,  I, -F) when "10101101001", 
		    to_sfixed(-0.895966,  I, -F) when "10101101010", 
		    to_sfixed(-0.897325,  I, -F) when "10101101011", 
		    to_sfixed(-0.898674,  I, -F) when "10101101100", 
		    to_sfixed(-0.900016,  I, -F) when "10101101101", 
		    to_sfixed(-0.901349,  I, -F) when "10101101110", 
		    to_sfixed(-0.902673,  I, -F) when "10101101111", 
		    to_sfixed(-0.903989,  I, -F) when "10101110000", 
		    to_sfixed(-0.905297,  I, -F) when "10101110001", 
		    to_sfixed(-0.906596,  I, -F) when "10101110010", 
		    to_sfixed(-0.907886,  I, -F) when "10101110011", 
		    to_sfixed(-0.909168,  I, -F) when "10101110100", 
		    to_sfixed(-0.910441,  I, -F) when "10101110101", 
		    to_sfixed(-0.911706,  I, -F) when "10101110110", 
		    to_sfixed(-0.912962,  I, -F) when "10101110111", 
		    to_sfixed(-0.914210,  I, -F) when "10101111000", 
		    to_sfixed(-0.915449,  I, -F) when "10101111001", 
		    to_sfixed(-0.916679,  I, -F) when "10101111010", 
		    to_sfixed(-0.917901,  I, -F) when "10101111011", 
		    to_sfixed(-0.919114,  I, -F) when "10101111100", 
		    to_sfixed(-0.920318,  I, -F) when "10101111101", 
		    to_sfixed(-0.921514,  I, -F) when "10101111110", 
		    to_sfixed(-0.922701,  I, -F) when "10101111111", 
		    to_sfixed(-0.923880,  I, -F) when "10110000000", 
		    to_sfixed(-0.925049,  I, -F) when "10110000001", 
		    to_sfixed(-0.926210,  I, -F) when "10110000010", 
		    to_sfixed(-0.927363,  I, -F) when "10110000011", 
		    to_sfixed(-0.928506,  I, -F) when "10110000100", 
		    to_sfixed(-0.929641,  I, -F) when "10110000101", 
		    to_sfixed(-0.930767,  I, -F) when "10110000110", 
		    to_sfixed(-0.931884,  I, -F) when "10110000111", 
		    to_sfixed(-0.932993,  I, -F) when "10110001000", 
		    to_sfixed(-0.934093,  I, -F) when "10110001001", 
		    to_sfixed(-0.935184,  I, -F) when "10110001010", 
		    to_sfixed(-0.936266,  I, -F) when "10110001011", 
		    to_sfixed(-0.937339,  I, -F) when "10110001100", 
		    to_sfixed(-0.938404,  I, -F) when "10110001101", 
		    to_sfixed(-0.939459,  I, -F) when "10110001110", 
		    to_sfixed(-0.940506,  I, -F) when "10110001111", 
		    to_sfixed(-0.941544,  I, -F) when "10110010000", 
		    to_sfixed(-0.942573,  I, -F) when "10110010001", 
		    to_sfixed(-0.943593,  I, -F) when "10110010010", 
		    to_sfixed(-0.944605,  I, -F) when "10110010011", 
		    to_sfixed(-0.945607,  I, -F) when "10110010100", 
		    to_sfixed(-0.946601,  I, -F) when "10110010101", 
		    to_sfixed(-0.947586,  I, -F) when "10110010110", 
		    to_sfixed(-0.948561,  I, -F) when "10110010111", 
		    to_sfixed(-0.949528,  I, -F) when "10110011000", 
		    to_sfixed(-0.950486,  I, -F) when "10110011001", 
		    to_sfixed(-0.951435,  I, -F) when "10110011010", 
		    to_sfixed(-0.952375,  I, -F) when "10110011011", 
		    to_sfixed(-0.953306,  I, -F) when "10110011100", 
		    to_sfixed(-0.954228,  I, -F) when "10110011101", 
		    to_sfixed(-0.955141,  I, -F) when "10110011110", 
		    to_sfixed(-0.956045,  I, -F) when "10110011111", 
		    to_sfixed(-0.956940,  I, -F) when "10110100000", 
		    to_sfixed(-0.957826,  I, -F) when "10110100001", 
		    to_sfixed(-0.958703,  I, -F) when "10110100010", 
		    to_sfixed(-0.959572,  I, -F) when "10110100011", 
		    to_sfixed(-0.960431,  I, -F) when "10110100100", 
		    to_sfixed(-0.961280,  I, -F) when "10110100101", 
		    to_sfixed(-0.962121,  I, -F) when "10110100110", 
		    to_sfixed(-0.962953,  I, -F) when "10110100111", 
		    to_sfixed(-0.963776,  I, -F) when "10110101000", 
		    to_sfixed(-0.964590,  I, -F) when "10110101001", 
		    to_sfixed(-0.965394,  I, -F) when "10110101010", 
		    to_sfixed(-0.966190,  I, -F) when "10110101011", 
		    to_sfixed(-0.966976,  I, -F) when "10110101100", 
		    to_sfixed(-0.967754,  I, -F) when "10110101101", 
		    to_sfixed(-0.968522,  I, -F) when "10110101110", 
		    to_sfixed(-0.969281,  I, -F) when "10110101111", 
		    to_sfixed(-0.970031,  I, -F) when "10110110000", 
		    to_sfixed(-0.970772,  I, -F) when "10110110001", 
		    to_sfixed(-0.971504,  I, -F) when "10110110010", 
		    to_sfixed(-0.972226,  I, -F) when "10110110011", 
		    to_sfixed(-0.972940,  I, -F) when "10110110100", 
		    to_sfixed(-0.973644,  I, -F) when "10110110101", 
		    to_sfixed(-0.974339,  I, -F) when "10110110110", 
		    to_sfixed(-0.975025,  I, -F) when "10110110111", 
		    to_sfixed(-0.975702,  I, -F) when "10110111000", 
		    to_sfixed(-0.976370,  I, -F) when "10110111001", 
		    to_sfixed(-0.977028,  I, -F) when "10110111010", 
		    to_sfixed(-0.977677,  I, -F) when "10110111011", 
		    to_sfixed(-0.978317,  I, -F) when "10110111100", 
		    to_sfixed(-0.978948,  I, -F) when "10110111101", 
		    to_sfixed(-0.979570,  I, -F) when "10110111110", 
		    to_sfixed(-0.980182,  I, -F) when "10110111111", 
		    to_sfixed(-0.980785,  I, -F) when "10111000000", 
		    to_sfixed(-0.981379,  I, -F) when "10111000001", 
		    to_sfixed(-0.981964,  I, -F) when "10111000010", 
		    to_sfixed(-0.982539,  I, -F) when "10111000011", 
		    to_sfixed(-0.983105,  I, -F) when "10111000100", 
		    to_sfixed(-0.983662,  I, -F) when "10111000101", 
		    to_sfixed(-0.984210,  I, -F) when "10111000110", 
		    to_sfixed(-0.984749,  I, -F) when "10111000111", 
		    to_sfixed(-0.985278,  I, -F) when "10111001000", 
		    to_sfixed(-0.985798,  I, -F) when "10111001001", 
		    to_sfixed(-0.986308,  I, -F) when "10111001010", 
		    to_sfixed(-0.986809,  I, -F) when "10111001011", 
		    to_sfixed(-0.987301,  I, -F) when "10111001100", 
		    to_sfixed(-0.987784,  I, -F) when "10111001101", 
		    to_sfixed(-0.988258,  I, -F) when "10111001110", 
		    to_sfixed(-0.988722,  I, -F) when "10111001111", 
		    to_sfixed(-0.989177,  I, -F) when "10111010000", 
		    to_sfixed(-0.989622,  I, -F) when "10111010001", 
		    to_sfixed(-0.990058,  I, -F) when "10111010010", 
		    to_sfixed(-0.990485,  I, -F) when "10111010011", 
		    to_sfixed(-0.990903,  I, -F) when "10111010100", 
		    to_sfixed(-0.991311,  I, -F) when "10111010101", 
		    to_sfixed(-0.991710,  I, -F) when "10111010110", 
		    to_sfixed(-0.992099,  I, -F) when "10111010111", 
		    to_sfixed(-0.992480,  I, -F) when "10111011000", 
		    to_sfixed(-0.992850,  I, -F) when "10111011001", 
		    to_sfixed(-0.993212,  I, -F) when "10111011010", 
		    to_sfixed(-0.993564,  I, -F) when "10111011011", 
		    to_sfixed(-0.993907,  I, -F) when "10111011100", 
		    to_sfixed(-0.994240,  I, -F) when "10111011101", 
		    to_sfixed(-0.994565,  I, -F) when "10111011110", 
		    to_sfixed(-0.994879,  I, -F) when "10111011111", 
		    to_sfixed(-0.995185,  I, -F) when "10111100000", 
		    to_sfixed(-0.995481,  I, -F) when "10111100001", 
		    to_sfixed(-0.995767,  I, -F) when "10111100010", 
		    to_sfixed(-0.996045,  I, -F) when "10111100011", 
		    to_sfixed(-0.996313,  I, -F) when "10111100100", 
		    to_sfixed(-0.996571,  I, -F) when "10111100101", 
		    to_sfixed(-0.996820,  I, -F) when "10111100110", 
		    to_sfixed(-0.997060,  I, -F) when "10111100111", 
		    to_sfixed(-0.997290,  I, -F) when "10111101000", 
		    to_sfixed(-0.997511,  I, -F) when "10111101001", 
		    to_sfixed(-0.997723,  I, -F) when "10111101010", 
		    to_sfixed(-0.997925,  I, -F) when "10111101011", 
		    to_sfixed(-0.998118,  I, -F) when "10111101100", 
		    to_sfixed(-0.998302,  I, -F) when "10111101101", 
		    to_sfixed(-0.998476,  I, -F) when "10111101110", 
		    to_sfixed(-0.998640,  I, -F) when "10111101111", 
		    to_sfixed(-0.998795,  I, -F) when "10111110000", 
		    to_sfixed(-0.998941,  I, -F) when "10111110001", 
		    to_sfixed(-0.999078,  I, -F) when "10111110010", 
		    to_sfixed(-0.999205,  I, -F) when "10111110011", 
		    to_sfixed(-0.999322,  I, -F) when "10111110100", 
		    to_sfixed(-0.999431,  I, -F) when "10111110101", 
		    to_sfixed(-0.999529,  I, -F) when "10111110110", 
		    to_sfixed(-0.999619,  I, -F) when "10111110111", 
		    to_sfixed(-0.999699,  I, -F) when "10111111000", 
		    to_sfixed(-0.999769,  I, -F) when "10111111001", 
		    to_sfixed(-0.999831,  I, -F) when "10111111010", 
		    to_sfixed(-0.999882,  I, -F) when "10111111011", 
		    to_sfixed(-0.999925,  I, -F) when "10111111100", 
		    to_sfixed(-0.999958,  I, -F) when "10111111101", 
		    to_sfixed(-0.999981,  I, -F) when "10111111110", 
		    to_sfixed(-0.999995,  I, -F) when "10111111111", 
		    to_sfixed(-1.000000,  I, -F) when "11000000000", 
		    to_sfixed(-0.999995,  I, -F) when "11000000001", 
		    to_sfixed(-0.999981,  I, -F) when "11000000010", 
		    to_sfixed(-0.999958,  I, -F) when "11000000011", 
		    to_sfixed(-0.999925,  I, -F) when "11000000100", 
		    to_sfixed(-0.999882,  I, -F) when "11000000101", 
		    to_sfixed(-0.999831,  I, -F) when "11000000110", 
		    to_sfixed(-0.999769,  I, -F) when "11000000111", 
		    to_sfixed(-0.999699,  I, -F) when "11000001000", 
		    to_sfixed(-0.999619,  I, -F) when "11000001001", 
		    to_sfixed(-0.999529,  I, -F) when "11000001010", 
		    to_sfixed(-0.999431,  I, -F) when "11000001011", 
		    to_sfixed(-0.999322,  I, -F) when "11000001100", 
		    to_sfixed(-0.999205,  I, -F) when "11000001101", 
		    to_sfixed(-0.999078,  I, -F) when "11000001110", 
		    to_sfixed(-0.998941,  I, -F) when "11000001111", 
		    to_sfixed(-0.998795,  I, -F) when "11000010000", 
		    to_sfixed(-0.998640,  I, -F) when "11000010001", 
		    to_sfixed(-0.998476,  I, -F) when "11000010010", 
		    to_sfixed(-0.998302,  I, -F) when "11000010011", 
		    to_sfixed(-0.998118,  I, -F) when "11000010100", 
		    to_sfixed(-0.997925,  I, -F) when "11000010101", 
		    to_sfixed(-0.997723,  I, -F) when "11000010110", 
		    to_sfixed(-0.997511,  I, -F) when "11000010111", 
		    to_sfixed(-0.997290,  I, -F) when "11000011000", 
		    to_sfixed(-0.997060,  I, -F) when "11000011001", 
		    to_sfixed(-0.996820,  I, -F) when "11000011010", 
		    to_sfixed(-0.996571,  I, -F) when "11000011011", 
		    to_sfixed(-0.996313,  I, -F) when "11000011100", 
		    to_sfixed(-0.996045,  I, -F) when "11000011101", 
		    to_sfixed(-0.995767,  I, -F) when "11000011110", 
		    to_sfixed(-0.995481,  I, -F) when "11000011111", 
		    to_sfixed(-0.995185,  I, -F) when "11000100000", 
		    to_sfixed(-0.994879,  I, -F) when "11000100001", 
		    to_sfixed(-0.994565,  I, -F) when "11000100010", 
		    to_sfixed(-0.994240,  I, -F) when "11000100011", 
		    to_sfixed(-0.993907,  I, -F) when "11000100100", 
		    to_sfixed(-0.993564,  I, -F) when "11000100101", 
		    to_sfixed(-0.993212,  I, -F) when "11000100110", 
		    to_sfixed(-0.992850,  I, -F) when "11000100111", 
		    to_sfixed(-0.992480,  I, -F) when "11000101000", 
		    to_sfixed(-0.992099,  I, -F) when "11000101001", 
		    to_sfixed(-0.991710,  I, -F) when "11000101010", 
		    to_sfixed(-0.991311,  I, -F) when "11000101011", 
		    to_sfixed(-0.990903,  I, -F) when "11000101100", 
		    to_sfixed(-0.990485,  I, -F) when "11000101101", 
		    to_sfixed(-0.990058,  I, -F) when "11000101110", 
		    to_sfixed(-0.989622,  I, -F) when "11000101111", 
		    to_sfixed(-0.989177,  I, -F) when "11000110000", 
		    to_sfixed(-0.988722,  I, -F) when "11000110001", 
		    to_sfixed(-0.988258,  I, -F) when "11000110010", 
		    to_sfixed(-0.987784,  I, -F) when "11000110011", 
		    to_sfixed(-0.987301,  I, -F) when "11000110100", 
		    to_sfixed(-0.986809,  I, -F) when "11000110101", 
		    to_sfixed(-0.986308,  I, -F) when "11000110110", 
		    to_sfixed(-0.985798,  I, -F) when "11000110111", 
		    to_sfixed(-0.985278,  I, -F) when "11000111000", 
		    to_sfixed(-0.984749,  I, -F) when "11000111001", 
		    to_sfixed(-0.984210,  I, -F) when "11000111010", 
		    to_sfixed(-0.983662,  I, -F) when "11000111011", 
		    to_sfixed(-0.983105,  I, -F) when "11000111100", 
		    to_sfixed(-0.982539,  I, -F) when "11000111101", 
		    to_sfixed(-0.981964,  I, -F) when "11000111110", 
		    to_sfixed(-0.981379,  I, -F) when "11000111111", 
		    to_sfixed(-0.980785,  I, -F) when "11001000000", 
		    to_sfixed(-0.980182,  I, -F) when "11001000001", 
		    to_sfixed(-0.979570,  I, -F) when "11001000010", 
		    to_sfixed(-0.978948,  I, -F) when "11001000011", 
		    to_sfixed(-0.978317,  I, -F) when "11001000100", 
		    to_sfixed(-0.977677,  I, -F) when "11001000101", 
		    to_sfixed(-0.977028,  I, -F) when "11001000110", 
		    to_sfixed(-0.976370,  I, -F) when "11001000111", 
		    to_sfixed(-0.975702,  I, -F) when "11001001000", 
		    to_sfixed(-0.975025,  I, -F) when "11001001001", 
		    to_sfixed(-0.974339,  I, -F) when "11001001010", 
		    to_sfixed(-0.973644,  I, -F) when "11001001011", 
		    to_sfixed(-0.972940,  I, -F) when "11001001100", 
		    to_sfixed(-0.972226,  I, -F) when "11001001101", 
		    to_sfixed(-0.971504,  I, -F) when "11001001110", 
		    to_sfixed(-0.970772,  I, -F) when "11001001111", 
		    to_sfixed(-0.970031,  I, -F) when "11001010000", 
		    to_sfixed(-0.969281,  I, -F) when "11001010001", 
		    to_sfixed(-0.968522,  I, -F) when "11001010010", 
		    to_sfixed(-0.967754,  I, -F) when "11001010011", 
		    to_sfixed(-0.966976,  I, -F) when "11001010100", 
		    to_sfixed(-0.966190,  I, -F) when "11001010101", 
		    to_sfixed(-0.965394,  I, -F) when "11001010110", 
		    to_sfixed(-0.964590,  I, -F) when "11001010111", 
		    to_sfixed(-0.963776,  I, -F) when "11001011000", 
		    to_sfixed(-0.962953,  I, -F) when "11001011001", 
		    to_sfixed(-0.962121,  I, -F) when "11001011010", 
		    to_sfixed(-0.961280,  I, -F) when "11001011011", 
		    to_sfixed(-0.960431,  I, -F) when "11001011100", 
		    to_sfixed(-0.959572,  I, -F) when "11001011101", 
		    to_sfixed(-0.958703,  I, -F) when "11001011110", 
		    to_sfixed(-0.957826,  I, -F) when "11001011111", 
		    to_sfixed(-0.956940,  I, -F) when "11001100000", 
		    to_sfixed(-0.956045,  I, -F) when "11001100001", 
		    to_sfixed(-0.955141,  I, -F) when "11001100010", 
		    to_sfixed(-0.954228,  I, -F) when "11001100011", 
		    to_sfixed(-0.953306,  I, -F) when "11001100100", 
		    to_sfixed(-0.952375,  I, -F) when "11001100101", 
		    to_sfixed(-0.951435,  I, -F) when "11001100110", 
		    to_sfixed(-0.950486,  I, -F) when "11001100111", 
		    to_sfixed(-0.949528,  I, -F) when "11001101000", 
		    to_sfixed(-0.948561,  I, -F) when "11001101001", 
		    to_sfixed(-0.947586,  I, -F) when "11001101010", 
		    to_sfixed(-0.946601,  I, -F) when "11001101011", 
		    to_sfixed(-0.945607,  I, -F) when "11001101100", 
		    to_sfixed(-0.944605,  I, -F) when "11001101101", 
		    to_sfixed(-0.943593,  I, -F) when "11001101110", 
		    to_sfixed(-0.942573,  I, -F) when "11001101111", 
		    to_sfixed(-0.941544,  I, -F) when "11001110000", 
		    to_sfixed(-0.940506,  I, -F) when "11001110001", 
		    to_sfixed(-0.939459,  I, -F) when "11001110010", 
		    to_sfixed(-0.938404,  I, -F) when "11001110011", 
		    to_sfixed(-0.937339,  I, -F) when "11001110100", 
		    to_sfixed(-0.936266,  I, -F) when "11001110101", 
		    to_sfixed(-0.935184,  I, -F) when "11001110110", 
		    to_sfixed(-0.934093,  I, -F) when "11001110111", 
		    to_sfixed(-0.932993,  I, -F) when "11001111000", 
		    to_sfixed(-0.931884,  I, -F) when "11001111001", 
		    to_sfixed(-0.930767,  I, -F) when "11001111010", 
		    to_sfixed(-0.929641,  I, -F) when "11001111011", 
		    to_sfixed(-0.928506,  I, -F) when "11001111100", 
		    to_sfixed(-0.927363,  I, -F) when "11001111101", 
		    to_sfixed(-0.926210,  I, -F) when "11001111110", 
		    to_sfixed(-0.925049,  I, -F) when "11001111111", 
		    to_sfixed(-0.923880,  I, -F) when "11010000000", 
		    to_sfixed(-0.922701,  I, -F) when "11010000001", 
		    to_sfixed(-0.921514,  I, -F) when "11010000010", 
		    to_sfixed(-0.920318,  I, -F) when "11010000011", 
		    to_sfixed(-0.919114,  I, -F) when "11010000100", 
		    to_sfixed(-0.917901,  I, -F) when "11010000101", 
		    to_sfixed(-0.916679,  I, -F) when "11010000110", 
		    to_sfixed(-0.915449,  I, -F) when "11010000111", 
		    to_sfixed(-0.914210,  I, -F) when "11010001000", 
		    to_sfixed(-0.912962,  I, -F) when "11010001001", 
		    to_sfixed(-0.911706,  I, -F) when "11010001010", 
		    to_sfixed(-0.910441,  I, -F) when "11010001011", 
		    to_sfixed(-0.909168,  I, -F) when "11010001100", 
		    to_sfixed(-0.907886,  I, -F) when "11010001101", 
		    to_sfixed(-0.906596,  I, -F) when "11010001110", 
		    to_sfixed(-0.905297,  I, -F) when "11010001111", 
		    to_sfixed(-0.903989,  I, -F) when "11010010000", 
		    to_sfixed(-0.902673,  I, -F) when "11010010001", 
		    to_sfixed(-0.901349,  I, -F) when "11010010010", 
		    to_sfixed(-0.900016,  I, -F) when "11010010011", 
		    to_sfixed(-0.898674,  I, -F) when "11010010100", 
		    to_sfixed(-0.897325,  I, -F) when "11010010101", 
		    to_sfixed(-0.895966,  I, -F) when "11010010110", 
		    to_sfixed(-0.894599,  I, -F) when "11010010111", 
		    to_sfixed(-0.893224,  I, -F) when "11010011000", 
		    to_sfixed(-0.891841,  I, -F) when "11010011001", 
		    to_sfixed(-0.890449,  I, -F) when "11010011010", 
		    to_sfixed(-0.889048,  I, -F) when "11010011011", 
		    to_sfixed(-0.887640,  I, -F) when "11010011100", 
		    to_sfixed(-0.886223,  I, -F) when "11010011101", 
		    to_sfixed(-0.884797,  I, -F) when "11010011110", 
		    to_sfixed(-0.883363,  I, -F) when "11010011111", 
		    to_sfixed(-0.881921,  I, -F) when "11010100000", 
		    to_sfixed(-0.880471,  I, -F) when "11010100001", 
		    to_sfixed(-0.879012,  I, -F) when "11010100010", 
		    to_sfixed(-0.877545,  I, -F) when "11010100011", 
		    to_sfixed(-0.876070,  I, -F) when "11010100100", 
		    to_sfixed(-0.874587,  I, -F) when "11010100101", 
		    to_sfixed(-0.873095,  I, -F) when "11010100110", 
		    to_sfixed(-0.871595,  I, -F) when "11010100111", 
		    to_sfixed(-0.870087,  I, -F) when "11010101000", 
		    to_sfixed(-0.868571,  I, -F) when "11010101001", 
		    to_sfixed(-0.867046,  I, -F) when "11010101010", 
		    to_sfixed(-0.865514,  I, -F) when "11010101011", 
		    to_sfixed(-0.863973,  I, -F) when "11010101100", 
		    to_sfixed(-0.862424,  I, -F) when "11010101101", 
		    to_sfixed(-0.860867,  I, -F) when "11010101110", 
		    to_sfixed(-0.859302,  I, -F) when "11010101111", 
		    to_sfixed(-0.857729,  I, -F) when "11010110000", 
		    to_sfixed(-0.856147,  I, -F) when "11010110001", 
		    to_sfixed(-0.854558,  I, -F) when "11010110010", 
		    to_sfixed(-0.852961,  I, -F) when "11010110011", 
		    to_sfixed(-0.851355,  I, -F) when "11010110100", 
		    to_sfixed(-0.849742,  I, -F) when "11010110101", 
		    to_sfixed(-0.848120,  I, -F) when "11010110110", 
		    to_sfixed(-0.846491,  I, -F) when "11010110111", 
		    to_sfixed(-0.844854,  I, -F) when "11010111000", 
		    to_sfixed(-0.843208,  I, -F) when "11010111001", 
		    to_sfixed(-0.841555,  I, -F) when "11010111010", 
		    to_sfixed(-0.839894,  I, -F) when "11010111011", 
		    to_sfixed(-0.838225,  I, -F) when "11010111100", 
		    to_sfixed(-0.836548,  I, -F) when "11010111101", 
		    to_sfixed(-0.834863,  I, -F) when "11010111110", 
		    to_sfixed(-0.833170,  I, -F) when "11010111111", 
		    to_sfixed(-0.831470,  I, -F) when "11011000000", 
		    to_sfixed(-0.829761,  I, -F) when "11011000001", 
		    to_sfixed(-0.828045,  I, -F) when "11011000010", 
		    to_sfixed(-0.826321,  I, -F) when "11011000011", 
		    to_sfixed(-0.824589,  I, -F) when "11011000100", 
		    to_sfixed(-0.822850,  I, -F) when "11011000101", 
		    to_sfixed(-0.821103,  I, -F) when "11011000110", 
		    to_sfixed(-0.819348,  I, -F) when "11011000111", 
		    to_sfixed(-0.817585,  I, -F) when "11011001000", 
		    to_sfixed(-0.815814,  I, -F) when "11011001001", 
		    to_sfixed(-0.814036,  I, -F) when "11011001010", 
		    to_sfixed(-0.812251,  I, -F) when "11011001011", 
		    to_sfixed(-0.810457,  I, -F) when "11011001100", 
		    to_sfixed(-0.808656,  I, -F) when "11011001101", 
		    to_sfixed(-0.806848,  I, -F) when "11011001110", 
		    to_sfixed(-0.805031,  I, -F) when "11011001111", 
		    to_sfixed(-0.803208,  I, -F) when "11011010000", 
		    to_sfixed(-0.801376,  I, -F) when "11011010001", 
		    to_sfixed(-0.799537,  I, -F) when "11011010010", 
		    to_sfixed(-0.797691,  I, -F) when "11011010011", 
		    to_sfixed(-0.795837,  I, -F) when "11011010100", 
		    to_sfixed(-0.793975,  I, -F) when "11011010101", 
		    to_sfixed(-0.792107,  I, -F) when "11011010110", 
		    to_sfixed(-0.790230,  I, -F) when "11011010111", 
		    to_sfixed(-0.788346,  I, -F) when "11011011000", 
		    to_sfixed(-0.786455,  I, -F) when "11011011001", 
		    to_sfixed(-0.784557,  I, -F) when "11011011010", 
		    to_sfixed(-0.782651,  I, -F) when "11011011011", 
		    to_sfixed(-0.780737,  I, -F) when "11011011100", 
		    to_sfixed(-0.778817,  I, -F) when "11011011101", 
		    to_sfixed(-0.776888,  I, -F) when "11011011110", 
		    to_sfixed(-0.774953,  I, -F) when "11011011111", 
		    to_sfixed(-0.773010,  I, -F) when "11011100000", 
		    to_sfixed(-0.771061,  I, -F) when "11011100001", 
		    to_sfixed(-0.769103,  I, -F) when "11011100010", 
		    to_sfixed(-0.767139,  I, -F) when "11011100011", 
		    to_sfixed(-0.765167,  I, -F) when "11011100100", 
		    to_sfixed(-0.763188,  I, -F) when "11011100101", 
		    to_sfixed(-0.761202,  I, -F) when "11011100110", 
		    to_sfixed(-0.759209,  I, -F) when "11011100111", 
		    to_sfixed(-0.757209,  I, -F) when "11011101000", 
		    to_sfixed(-0.755201,  I, -F) when "11011101001", 
		    to_sfixed(-0.753187,  I, -F) when "11011101010", 
		    to_sfixed(-0.751165,  I, -F) when "11011101011", 
		    to_sfixed(-0.749136,  I, -F) when "11011101100", 
		    to_sfixed(-0.747101,  I, -F) when "11011101101", 
		    to_sfixed(-0.745058,  I, -F) when "11011101110", 
		    to_sfixed(-0.743008,  I, -F) when "11011101111", 
		    to_sfixed(-0.740951,  I, -F) when "11011110000", 
		    to_sfixed(-0.738887,  I, -F) when "11011110001", 
		    to_sfixed(-0.736817,  I, -F) when "11011110010", 
		    to_sfixed(-0.734739,  I, -F) when "11011110011", 
		    to_sfixed(-0.732654,  I, -F) when "11011110100", 
		    to_sfixed(-0.730563,  I, -F) when "11011110101", 
		    to_sfixed(-0.728464,  I, -F) when "11011110110", 
		    to_sfixed(-0.726359,  I, -F) when "11011110111", 
		    to_sfixed(-0.724247,  I, -F) when "11011111000", 
		    to_sfixed(-0.722128,  I, -F) when "11011111001", 
		    to_sfixed(-0.720003,  I, -F) when "11011111010", 
		    to_sfixed(-0.717870,  I, -F) when "11011111011", 
		    to_sfixed(-0.715731,  I, -F) when "11011111100", 
		    to_sfixed(-0.713585,  I, -F) when "11011111101", 
		    to_sfixed(-0.711432,  I, -F) when "11011111110", 
		    to_sfixed(-0.709273,  I, -F) when "11011111111", 
		    to_sfixed(-0.707107,  I, -F) when "11100000000", 
		    to_sfixed(-0.704934,  I, -F) when "11100000001", 
		    to_sfixed(-0.702755,  I, -F) when "11100000010", 
		    to_sfixed(-0.700569,  I, -F) when "11100000011", 
		    to_sfixed(-0.698376,  I, -F) when "11100000100", 
		    to_sfixed(-0.696177,  I, -F) when "11100000101", 
		    to_sfixed(-0.693971,  I, -F) when "11100000110", 
		    to_sfixed(-0.691759,  I, -F) when "11100000111", 
		    to_sfixed(-0.689541,  I, -F) when "11100001000", 
		    to_sfixed(-0.687315,  I, -F) when "11100001001", 
		    to_sfixed(-0.685084,  I, -F) when "11100001010", 
		    to_sfixed(-0.682846,  I, -F) when "11100001011", 
		    to_sfixed(-0.680601,  I, -F) when "11100001100", 
		    to_sfixed(-0.678350,  I, -F) when "11100001101", 
		    to_sfixed(-0.676093,  I, -F) when "11100001110", 
		    to_sfixed(-0.673829,  I, -F) when "11100001111", 
		    to_sfixed(-0.671559,  I, -F) when "11100010000", 
		    to_sfixed(-0.669283,  I, -F) when "11100010001", 
		    to_sfixed(-0.667000,  I, -F) when "11100010010", 
		    to_sfixed(-0.664711,  I, -F) when "11100010011", 
		    to_sfixed(-0.662416,  I, -F) when "11100010100", 
		    to_sfixed(-0.660114,  I, -F) when "11100010101", 
		    to_sfixed(-0.657807,  I, -F) when "11100010110", 
		    to_sfixed(-0.655493,  I, -F) when "11100010111", 
		    to_sfixed(-0.653173,  I, -F) when "11100011000", 
		    to_sfixed(-0.650847,  I, -F) when "11100011001", 
		    to_sfixed(-0.648514,  I, -F) when "11100011010", 
		    to_sfixed(-0.646176,  I, -F) when "11100011011", 
		    to_sfixed(-0.643832,  I, -F) when "11100011100", 
		    to_sfixed(-0.641481,  I, -F) when "11100011101", 
		    to_sfixed(-0.639124,  I, -F) when "11100011110", 
		    to_sfixed(-0.636762,  I, -F) when "11100011111", 
		    to_sfixed(-0.634393,  I, -F) when "11100100000", 
		    to_sfixed(-0.632019,  I, -F) when "11100100001", 
		    to_sfixed(-0.629638,  I, -F) when "11100100010", 
		    to_sfixed(-0.627252,  I, -F) when "11100100011", 
		    to_sfixed(-0.624859,  I, -F) when "11100100100", 
		    to_sfixed(-0.622461,  I, -F) when "11100100101", 
		    to_sfixed(-0.620057,  I, -F) when "11100100110", 
		    to_sfixed(-0.617647,  I, -F) when "11100100111", 
		    to_sfixed(-0.615232,  I, -F) when "11100101000", 
		    to_sfixed(-0.612810,  I, -F) when "11100101001", 
		    to_sfixed(-0.610383,  I, -F) when "11100101010", 
		    to_sfixed(-0.607950,  I, -F) when "11100101011", 
		    to_sfixed(-0.605511,  I, -F) when "11100101100", 
		    to_sfixed(-0.603067,  I, -F) when "11100101101", 
		    to_sfixed(-0.600616,  I, -F) when "11100101110", 
		    to_sfixed(-0.598161,  I, -F) when "11100101111", 
		    to_sfixed(-0.595699,  I, -F) when "11100110000", 
		    to_sfixed(-0.593232,  I, -F) when "11100110001", 
		    to_sfixed(-0.590760,  I, -F) when "11100110010", 
		    to_sfixed(-0.588282,  I, -F) when "11100110011", 
		    to_sfixed(-0.585798,  I, -F) when "11100110100", 
		    to_sfixed(-0.583309,  I, -F) when "11100110101", 
		    to_sfixed(-0.580814,  I, -F) when "11100110110", 
		    to_sfixed(-0.578314,  I, -F) when "11100110111", 
		    to_sfixed(-0.575808,  I, -F) when "11100111000", 
		    to_sfixed(-0.573297,  I, -F) when "11100111001", 
		    to_sfixed(-0.570781,  I, -F) when "11100111010", 
		    to_sfixed(-0.568259,  I, -F) when "11100111011", 
		    to_sfixed(-0.565732,  I, -F) when "11100111100", 
		    to_sfixed(-0.563199,  I, -F) when "11100111101", 
		    to_sfixed(-0.560662,  I, -F) when "11100111110", 
		    to_sfixed(-0.558119,  I, -F) when "11100111111", 
		    to_sfixed(-0.555570,  I, -F) when "11101000000", 
		    to_sfixed(-0.553017,  I, -F) when "11101000001", 
		    to_sfixed(-0.550458,  I, -F) when "11101000010", 
		    to_sfixed(-0.547894,  I, -F) when "11101000011", 
		    to_sfixed(-0.545325,  I, -F) when "11101000100", 
		    to_sfixed(-0.542751,  I, -F) when "11101000101", 
		    to_sfixed(-0.540171,  I, -F) when "11101000110", 
		    to_sfixed(-0.537587,  I, -F) when "11101000111", 
		    to_sfixed(-0.534998,  I, -F) when "11101001000", 
		    to_sfixed(-0.532403,  I, -F) when "11101001001", 
		    to_sfixed(-0.529804,  I, -F) when "11101001010", 
		    to_sfixed(-0.527199,  I, -F) when "11101001011", 
		    to_sfixed(-0.524590,  I, -F) when "11101001100", 
		    to_sfixed(-0.521975,  I, -F) when "11101001101", 
		    to_sfixed(-0.519356,  I, -F) when "11101001110", 
		    to_sfixed(-0.516732,  I, -F) when "11101001111", 
		    to_sfixed(-0.514103,  I, -F) when "11101010000", 
		    to_sfixed(-0.511469,  I, -F) when "11101010001", 
		    to_sfixed(-0.508830,  I, -F) when "11101010010", 
		    to_sfixed(-0.506187,  I, -F) when "11101010011", 
		    to_sfixed(-0.503538,  I, -F) when "11101010100", 
		    to_sfixed(-0.500885,  I, -F) when "11101010101", 
		    to_sfixed(-0.498228,  I, -F) when "11101010110", 
		    to_sfixed(-0.495565,  I, -F) when "11101010111", 
		    to_sfixed(-0.492898,  I, -F) when "11101011000", 
		    to_sfixed(-0.490226,  I, -F) when "11101011001", 
		    to_sfixed(-0.487550,  I, -F) when "11101011010", 
		    to_sfixed(-0.484869,  I, -F) when "11101011011", 
		    to_sfixed(-0.482184,  I, -F) when "11101011100", 
		    to_sfixed(-0.479494,  I, -F) when "11101011101", 
		    to_sfixed(-0.476799,  I, -F) when "11101011110", 
		    to_sfixed(-0.474100,  I, -F) when "11101011111", 
		    to_sfixed(-0.471397,  I, -F) when "11101100000", 
		    to_sfixed(-0.468689,  I, -F) when "11101100001", 
		    to_sfixed(-0.465976,  I, -F) when "11101100010", 
		    to_sfixed(-0.463260,  I, -F) when "11101100011", 
		    to_sfixed(-0.460539,  I, -F) when "11101100100", 
		    to_sfixed(-0.457813,  I, -F) when "11101100101", 
		    to_sfixed(-0.455084,  I, -F) when "11101100110", 
		    to_sfixed(-0.452350,  I, -F) when "11101100111", 
		    to_sfixed(-0.449611,  I, -F) when "11101101000", 
		    to_sfixed(-0.446869,  I, -F) when "11101101001", 
		    to_sfixed(-0.444122,  I, -F) when "11101101010", 
		    to_sfixed(-0.441371,  I, -F) when "11101101011", 
		    to_sfixed(-0.438616,  I, -F) when "11101101100", 
		    to_sfixed(-0.435857,  I, -F) when "11101101101", 
		    to_sfixed(-0.433094,  I, -F) when "11101101110", 
		    to_sfixed(-0.430326,  I, -F) when "11101101111", 
		    to_sfixed(-0.427555,  I, -F) when "11101110000", 
		    to_sfixed(-0.424780,  I, -F) when "11101110001", 
		    to_sfixed(-0.422000,  I, -F) when "11101110010", 
		    to_sfixed(-0.419217,  I, -F) when "11101110011", 
		    to_sfixed(-0.416430,  I, -F) when "11101110100", 
		    to_sfixed(-0.413638,  I, -F) when "11101110101", 
		    to_sfixed(-0.410843,  I, -F) when "11101110110", 
		    to_sfixed(-0.408044,  I, -F) when "11101110111", 
		    to_sfixed(-0.405241,  I, -F) when "11101111000", 
		    to_sfixed(-0.402435,  I, -F) when "11101111001", 
		    to_sfixed(-0.399624,  I, -F) when "11101111010", 
		    to_sfixed(-0.396810,  I, -F) when "11101111011", 
		    to_sfixed(-0.393992,  I, -F) when "11101111100", 
		    to_sfixed(-0.391170,  I, -F) when "11101111101", 
		    to_sfixed(-0.388345,  I, -F) when "11101111110", 
		    to_sfixed(-0.385516,  I, -F) when "11101111111", 
		    to_sfixed(-0.382683,  I, -F) when "11110000000", 
		    to_sfixed(-0.379847,  I, -F) when "11110000001", 
		    to_sfixed(-0.377007,  I, -F) when "11110000010", 
		    to_sfixed(-0.374164,  I, -F) when "11110000011", 
		    to_sfixed(-0.371317,  I, -F) when "11110000100", 
		    to_sfixed(-0.368467,  I, -F) when "11110000101", 
		    to_sfixed(-0.365613,  I, -F) when "11110000110", 
		    to_sfixed(-0.362756,  I, -F) when "11110000111", 
		    to_sfixed(-0.359895,  I, -F) when "11110001000", 
		    to_sfixed(-0.357031,  I, -F) when "11110001001", 
		    to_sfixed(-0.354164,  I, -F) when "11110001010", 
		    to_sfixed(-0.351293,  I, -F) when "11110001011", 
		    to_sfixed(-0.348419,  I, -F) when "11110001100", 
		    to_sfixed(-0.345541,  I, -F) when "11110001101", 
		    to_sfixed(-0.342661,  I, -F) when "11110001110", 
		    to_sfixed(-0.339777,  I, -F) when "11110001111", 
		    to_sfixed(-0.336890,  I, -F) when "11110010000", 
		    to_sfixed(-0.334000,  I, -F) when "11110010001", 
		    to_sfixed(-0.331106,  I, -F) when "11110010010", 
		    to_sfixed(-0.328210,  I, -F) when "11110010011", 
		    to_sfixed(-0.325310,  I, -F) when "11110010100", 
		    to_sfixed(-0.322408,  I, -F) when "11110010101", 
		    to_sfixed(-0.319502,  I, -F) when "11110010110", 
		    to_sfixed(-0.316593,  I, -F) when "11110010111", 
		    to_sfixed(-0.313682,  I, -F) when "11110011000", 
		    to_sfixed(-0.310767,  I, -F) when "11110011001", 
		    to_sfixed(-0.307850,  I, -F) when "11110011010", 
		    to_sfixed(-0.304929,  I, -F) when "11110011011", 
		    to_sfixed(-0.302006,  I, -F) when "11110011100", 
		    to_sfixed(-0.299080,  I, -F) when "11110011101", 
		    to_sfixed(-0.296151,  I, -F) when "11110011110", 
		    to_sfixed(-0.293219,  I, -F) when "11110011111", 
		    to_sfixed(-0.290285,  I, -F) when "11110100000", 
		    to_sfixed(-0.287347,  I, -F) when "11110100001", 
		    to_sfixed(-0.284408,  I, -F) when "11110100010", 
		    to_sfixed(-0.281465,  I, -F) when "11110100011", 
		    to_sfixed(-0.278520,  I, -F) when "11110100100", 
		    to_sfixed(-0.275572,  I, -F) when "11110100101", 
		    to_sfixed(-0.272621,  I, -F) when "11110100110", 
		    to_sfixed(-0.269668,  I, -F) when "11110100111", 
		    to_sfixed(-0.266713,  I, -F) when "11110101000", 
		    to_sfixed(-0.263755,  I, -F) when "11110101001", 
		    to_sfixed(-0.260794,  I, -F) when "11110101010", 
		    to_sfixed(-0.257831,  I, -F) when "11110101011", 
		    to_sfixed(-0.254866,  I, -F) when "11110101100", 
		    to_sfixed(-0.251898,  I, -F) when "11110101101", 
		    to_sfixed(-0.248928,  I, -F) when "11110101110", 
		    to_sfixed(-0.245955,  I, -F) when "11110101111", 
		    to_sfixed(-0.242980,  I, -F) when "11110110000", 
		    to_sfixed(-0.240003,  I, -F) when "11110110001", 
		    to_sfixed(-0.237024,  I, -F) when "11110110010", 
		    to_sfixed(-0.234042,  I, -F) when "11110110011", 
		    to_sfixed(-0.231058,  I, -F) when "11110110100", 
		    to_sfixed(-0.228072,  I, -F) when "11110110101", 
		    to_sfixed(-0.225084,  I, -F) when "11110110110", 
		    to_sfixed(-0.222094,  I, -F) when "11110110111", 
		    to_sfixed(-0.219101,  I, -F) when "11110111000", 
		    to_sfixed(-0.216107,  I, -F) when "11110111001", 
		    to_sfixed(-0.213110,  I, -F) when "11110111010", 
		    to_sfixed(-0.210112,  I, -F) when "11110111011", 
		    to_sfixed(-0.207111,  I, -F) when "11110111100", 
		    to_sfixed(-0.204109,  I, -F) when "11110111101", 
		    to_sfixed(-0.201105,  I, -F) when "11110111110", 
		    to_sfixed(-0.198098,  I, -F) when "11110111111", 
		    to_sfixed(-0.195090,  I, -F) when "11111000000", 
		    to_sfixed(-0.192080,  I, -F) when "11111000001", 
		    to_sfixed(-0.189069,  I, -F) when "11111000010", 
		    to_sfixed(-0.186055,  I, -F) when "11111000011", 
		    to_sfixed(-0.183040,  I, -F) when "11111000100", 
		    to_sfixed(-0.180023,  I, -F) when "11111000101", 
		    to_sfixed(-0.177004,  I, -F) when "11111000110", 
		    to_sfixed(-0.173984,  I, -F) when "11111000111", 
		    to_sfixed(-0.170962,  I, -F) when "11111001000", 
		    to_sfixed(-0.167938,  I, -F) when "11111001001", 
		    to_sfixed(-0.164913,  I, -F) when "11111001010", 
		    to_sfixed(-0.161886,  I, -F) when "11111001011", 
		    to_sfixed(-0.158858,  I, -F) when "11111001100", 
		    to_sfixed(-0.155828,  I, -F) when "11111001101", 
		    to_sfixed(-0.152797,  I, -F) when "11111001110", 
		    to_sfixed(-0.149765,  I, -F) when "11111001111", 
		    to_sfixed(-0.146730,  I, -F) when "11111010000", 
		    to_sfixed(-0.143695,  I, -F) when "11111010001", 
		    to_sfixed(-0.140658,  I, -F) when "11111010010", 
		    to_sfixed(-0.137620,  I, -F) when "11111010011", 
		    to_sfixed(-0.134581,  I, -F) when "11111010100", 
		    to_sfixed(-0.131540,  I, -F) when "11111010101", 
		    to_sfixed(-0.128498,  I, -F) when "11111010110", 
		    to_sfixed(-0.125455,  I, -F) when "11111010111", 
		    to_sfixed(-0.122411,  I, -F) when "11111011000", 
		    to_sfixed(-0.119365,  I, -F) when "11111011001", 
		    to_sfixed(-0.116319,  I, -F) when "11111011010", 
		    to_sfixed(-0.113271,  I, -F) when "11111011011", 
		    to_sfixed(-0.110222,  I, -F) when "11111011100", 
		    to_sfixed(-0.107172,  I, -F) when "11111011101", 
		    to_sfixed(-0.104122,  I, -F) when "11111011110", 
		    to_sfixed(-0.101070,  I, -F) when "11111011111", 
		    to_sfixed(-0.098017,  I, -F) when "11111100000", 
		    to_sfixed(-0.094963,  I, -F) when "11111100001", 
		    to_sfixed(-0.091909,  I, -F) when "11111100010", 
		    to_sfixed(-0.088854,  I, -F) when "11111100011", 
		    to_sfixed(-0.085797,  I, -F) when "11111100100", 
		    to_sfixed(-0.082740,  I, -F) when "11111100101", 
		    to_sfixed(-0.079682,  I, -F) when "11111100110", 
		    to_sfixed(-0.076624,  I, -F) when "11111100111", 
		    to_sfixed(-0.073565,  I, -F) when "11111101000", 
		    to_sfixed(-0.070505,  I, -F) when "11111101001", 
		    to_sfixed(-0.067444,  I, -F) when "11111101010", 
		    to_sfixed(-0.064383,  I, -F) when "11111101011", 
		    to_sfixed(-0.061321,  I, -F) when "11111101100", 
		    to_sfixed(-0.058258,  I, -F) when "11111101101", 
		    to_sfixed(-0.055195,  I, -F) when "11111101110", 
		    to_sfixed(-0.052132,  I, -F) when "11111101111", 
		    to_sfixed(-0.049068,  I, -F) when "11111110000", 
		    to_sfixed(-0.046003,  I, -F) when "11111110001", 
		    to_sfixed(-0.042938,  I, -F) when "11111110010", 
		    to_sfixed(-0.039873,  I, -F) when "11111110011", 
		    to_sfixed(-0.036807,  I, -F) when "11111110100", 
		    to_sfixed(-0.033741,  I, -F) when "11111110101", 
		    to_sfixed(-0.030675,  I, -F) when "11111110110", 
		    to_sfixed(-0.027608,  I, -F) when "11111110111", 
		    to_sfixed(-0.024541,  I, -F) when "11111111000", 
		    to_sfixed(-0.021474,  I, -F) when "11111111001", 
		    to_sfixed(-0.018407,  I, -F) when "11111111010", 
		    to_sfixed(-0.015339,  I, -F) when "11111111011", 
		    to_sfixed(-0.012272,  I, -F) when "11111111100", 
		    to_sfixed(-0.009204,  I, -F) when "11111111101", 
		    to_sfixed(-0.006136,  I, -F) when "11111111110", 
		    to_sfixed(-0.003068,  I, -F) when "11111111111", 
		    to_sfixed(0, I, -F) when others;
    
end architecture tabela_sin;

