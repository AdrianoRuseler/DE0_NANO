library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;


entity tabela_sin is
    generic (-- constant THETA_MAX : integer := 380808000;  --eqquivalente a 2*pi
                 constant n_bits_phase : integer :=16;  --numero de bits que representa a fase da rede
                 constant n_bits_c: integer := 16  --numero de bits da portadora    
             );
    port (clk : in std_logic;
          theta: in std_logic_vector(n_bits_phase-1 downto 0);
          va : out std_logic_vector(n_bits_c-1 downto 0)
          );
end tabela_sin;

architecture tabela_sin of tabela_sin is
    signal id : std_logic_vector(10 downto 0);
    signal sin : std_logic_vector(n_bits_c-1 downto 0);
	 signal va_int : std_logic_vector(n_bits_c*2-1 downto 0);
begin 
    
  id <= theta(n_bits_phase-1 downto n_bits_phase-11); -- 15 downto 5 - resolução do pwm?
   -- id <= theta; 
    
    process(clk)
    begin
        if rising_edge(clk) then
				va <= sin;
        end if;
    end process;
with id select
  sin <= 		    std_logic_vector(to_unsigned(668, n_bits_c)) when "00000000000", 
		    std_logic_vector(to_unsigned(669, n_bits_c)) when "00000000001", 
		    std_logic_vector(to_unsigned(671, n_bits_c)) when "00000000010", 
		    std_logic_vector(to_unsigned(672, n_bits_c)) when "00000000011", 
		    std_logic_vector(to_unsigned(674, n_bits_c)) when "00000000100", 
		    std_logic_vector(to_unsigned(676, n_bits_c)) when "00000000101", 
		    std_logic_vector(to_unsigned(677, n_bits_c)) when "00000000110", 
		    std_logic_vector(to_unsigned(679, n_bits_c)) when "00000000111", 
		    std_logic_vector(to_unsigned(681, n_bits_c)) when "00000001000", 
		    std_logic_vector(to_unsigned(682, n_bits_c)) when "00000001001", 
		    std_logic_vector(to_unsigned(684, n_bits_c)) when "00000001010", 
		    std_logic_vector(to_unsigned(686, n_bits_c)) when "00000001011", 
		    std_logic_vector(to_unsigned(687, n_bits_c)) when "00000001100", 
		    std_logic_vector(to_unsigned(689, n_bits_c)) when "00000001101", 
		    std_logic_vector(to_unsigned(691, n_bits_c)) when "00000001110", 
		    std_logic_vector(to_unsigned(692, n_bits_c)) when "00000001111", 
		    std_logic_vector(to_unsigned(694, n_bits_c)) when "00000010000", 
		    std_logic_vector(to_unsigned(696, n_bits_c)) when "00000010001", 
		    std_logic_vector(to_unsigned(697, n_bits_c)) when "00000010010", 
		    std_logic_vector(to_unsigned(699, n_bits_c)) when "00000010011", 
		    std_logic_vector(to_unsigned(701, n_bits_c)) when "00000010100", 
		    std_logic_vector(to_unsigned(702, n_bits_c)) when "00000010101", 
		    std_logic_vector(to_unsigned(704, n_bits_c)) when "00000010110", 
		    std_logic_vector(to_unsigned(706, n_bits_c)) when "00000010111", 
		    std_logic_vector(to_unsigned(707, n_bits_c)) when "00000011000", 
		    std_logic_vector(to_unsigned(709, n_bits_c)) when "00000011001", 
		    std_logic_vector(to_unsigned(711, n_bits_c)) when "00000011010", 
		    std_logic_vector(to_unsigned(712, n_bits_c)) when "00000011011", 
		    std_logic_vector(to_unsigned(714, n_bits_c)) when "00000011100", 
		    std_logic_vector(to_unsigned(716, n_bits_c)) when "00000011101", 
		    std_logic_vector(to_unsigned(717, n_bits_c)) when "00000011110", 
		    std_logic_vector(to_unsigned(719, n_bits_c)) when "00000011111", 
		    std_logic_vector(to_unsigned(721, n_bits_c)) when "00000100000", 
		    std_logic_vector(to_unsigned(722, n_bits_c)) when "00000100001", 
		    std_logic_vector(to_unsigned(724, n_bits_c)) when "00000100010", 
		    std_logic_vector(to_unsigned(726, n_bits_c)) when "00000100011", 
		    std_logic_vector(to_unsigned(727, n_bits_c)) when "00000100100", 
		    std_logic_vector(to_unsigned(729, n_bits_c)) when "00000100101", 
		    std_logic_vector(to_unsigned(731, n_bits_c)) when "00000100110", 
		    std_logic_vector(to_unsigned(732, n_bits_c)) when "00000100111", 
		    std_logic_vector(to_unsigned(734, n_bits_c)) when "00000101000", 
		    std_logic_vector(to_unsigned(736, n_bits_c)) when "00000101001", 
		    std_logic_vector(to_unsigned(737, n_bits_c)) when "00000101010", 
		    std_logic_vector(to_unsigned(739, n_bits_c)) when "00000101011", 
		    std_logic_vector(to_unsigned(741, n_bits_c)) when "00000101100", 
		    std_logic_vector(to_unsigned(742, n_bits_c)) when "00000101101", 
		    std_logic_vector(to_unsigned(744, n_bits_c)) when "00000101110", 
		    std_logic_vector(to_unsigned(746, n_bits_c)) when "00000101111", 
		    std_logic_vector(to_unsigned(747, n_bits_c)) when "00000110000", 
		    std_logic_vector(to_unsigned(749, n_bits_c)) when "00000110001", 
		    std_logic_vector(to_unsigned(750, n_bits_c)) when "00000110010", 
		    std_logic_vector(to_unsigned(752, n_bits_c)) when "00000110011", 
		    std_logic_vector(to_unsigned(754, n_bits_c)) when "00000110100", 
		    std_logic_vector(to_unsigned(755, n_bits_c)) when "00000110101", 
		    std_logic_vector(to_unsigned(757, n_bits_c)) when "00000110110", 
		    std_logic_vector(to_unsigned(759, n_bits_c)) when "00000110111", 
		    std_logic_vector(to_unsigned(760, n_bits_c)) when "00000111000", 
		    std_logic_vector(to_unsigned(762, n_bits_c)) when "00000111001", 
		    std_logic_vector(to_unsigned(764, n_bits_c)) when "00000111010", 
		    std_logic_vector(to_unsigned(765, n_bits_c)) when "00000111011", 
		    std_logic_vector(to_unsigned(767, n_bits_c)) when "00000111100", 
		    std_logic_vector(to_unsigned(769, n_bits_c)) when "00000111101", 
		    std_logic_vector(to_unsigned(770, n_bits_c)) when "00000111110", 
		    std_logic_vector(to_unsigned(772, n_bits_c)) when "00000111111", 
		    std_logic_vector(to_unsigned(773, n_bits_c)) when "00001000000", 
		    std_logic_vector(to_unsigned(775, n_bits_c)) when "00001000001", 
		    std_logic_vector(to_unsigned(777, n_bits_c)) when "00001000010", 
		    std_logic_vector(to_unsigned(778, n_bits_c)) when "00001000011", 
		    std_logic_vector(to_unsigned(780, n_bits_c)) when "00001000100", 
		    std_logic_vector(to_unsigned(782, n_bits_c)) when "00001000101", 
		    std_logic_vector(to_unsigned(783, n_bits_c)) when "00001000110", 
		    std_logic_vector(to_unsigned(785, n_bits_c)) when "00001000111", 
		    std_logic_vector(to_unsigned(787, n_bits_c)) when "00001001000", 
		    std_logic_vector(to_unsigned(788, n_bits_c)) when "00001001001", 
		    std_logic_vector(to_unsigned(790, n_bits_c)) when "00001001010", 
		    std_logic_vector(to_unsigned(791, n_bits_c)) when "00001001011", 
		    std_logic_vector(to_unsigned(793, n_bits_c)) when "00001001100", 
		    std_logic_vector(to_unsigned(795, n_bits_c)) when "00001001101", 
		    std_logic_vector(to_unsigned(796, n_bits_c)) when "00001001110", 
		    std_logic_vector(to_unsigned(798, n_bits_c)) when "00001001111", 
		    std_logic_vector(to_unsigned(799, n_bits_c)) when "00001010000", 
		    std_logic_vector(to_unsigned(801, n_bits_c)) when "00001010001", 
		    std_logic_vector(to_unsigned(803, n_bits_c)) when "00001010010", 
		    std_logic_vector(to_unsigned(804, n_bits_c)) when "00001010011", 
		    std_logic_vector(to_unsigned(806, n_bits_c)) when "00001010100", 
		    std_logic_vector(to_unsigned(808, n_bits_c)) when "00001010101", 
		    std_logic_vector(to_unsigned(809, n_bits_c)) when "00001010110", 
		    std_logic_vector(to_unsigned(811, n_bits_c)) when "00001010111", 
		    std_logic_vector(to_unsigned(812, n_bits_c)) when "00001011000", 
		    std_logic_vector(to_unsigned(814, n_bits_c)) when "00001011001", 
		    std_logic_vector(to_unsigned(816, n_bits_c)) when "00001011010", 
		    std_logic_vector(to_unsigned(817, n_bits_c)) when "00001011011", 
		    std_logic_vector(to_unsigned(819, n_bits_c)) when "00001011100", 
		    std_logic_vector(to_unsigned(820, n_bits_c)) when "00001011101", 
		    std_logic_vector(to_unsigned(822, n_bits_c)) when "00001011110", 
		    std_logic_vector(to_unsigned(824, n_bits_c)) when "00001011111", 
		    std_logic_vector(to_unsigned(825, n_bits_c)) when "00001100000", 
		    std_logic_vector(to_unsigned(827, n_bits_c)) when "00001100001", 
		    std_logic_vector(to_unsigned(828, n_bits_c)) when "00001100010", 
		    std_logic_vector(to_unsigned(830, n_bits_c)) when "00001100011", 
		    std_logic_vector(to_unsigned(832, n_bits_c)) when "00001100100", 
		    std_logic_vector(to_unsigned(833, n_bits_c)) when "00001100101", 
		    std_logic_vector(to_unsigned(835, n_bits_c)) when "00001100110", 
		    std_logic_vector(to_unsigned(836, n_bits_c)) when "00001100111", 
		    std_logic_vector(to_unsigned(838, n_bits_c)) when "00001101000", 
		    std_logic_vector(to_unsigned(839, n_bits_c)) when "00001101001", 
		    std_logic_vector(to_unsigned(841, n_bits_c)) when "00001101010", 
		    std_logic_vector(to_unsigned(843, n_bits_c)) when "00001101011", 
		    std_logic_vector(to_unsigned(844, n_bits_c)) when "00001101100", 
		    std_logic_vector(to_unsigned(846, n_bits_c)) when "00001101101", 
		    std_logic_vector(to_unsigned(847, n_bits_c)) when "00001101110", 
		    std_logic_vector(to_unsigned(849, n_bits_c)) when "00001101111", 
		    std_logic_vector(to_unsigned(850, n_bits_c)) when "00001110000", 
		    std_logic_vector(to_unsigned(852, n_bits_c)) when "00001110001", 
		    std_logic_vector(to_unsigned(854, n_bits_c)) when "00001110010", 
		    std_logic_vector(to_unsigned(855, n_bits_c)) when "00001110011", 
		    std_logic_vector(to_unsigned(857, n_bits_c)) when "00001110100", 
		    std_logic_vector(to_unsigned(858, n_bits_c)) when "00001110101", 
		    std_logic_vector(to_unsigned(860, n_bits_c)) when "00001110110", 
		    std_logic_vector(to_unsigned(861, n_bits_c)) when "00001110111", 
		    std_logic_vector(to_unsigned(863, n_bits_c)) when "00001111000", 
		    std_logic_vector(to_unsigned(865, n_bits_c)) when "00001111001", 
		    std_logic_vector(to_unsigned(866, n_bits_c)) when "00001111010", 
		    std_logic_vector(to_unsigned(868, n_bits_c)) when "00001111011", 
		    std_logic_vector(to_unsigned(869, n_bits_c)) when "00001111100", 
		    std_logic_vector(to_unsigned(871, n_bits_c)) when "00001111101", 
		    std_logic_vector(to_unsigned(872, n_bits_c)) when "00001111110", 
		    std_logic_vector(to_unsigned(874, n_bits_c)) when "00001111111", 
		    std_logic_vector(to_unsigned(875, n_bits_c)) when "00010000000", 
		    std_logic_vector(to_unsigned(877, n_bits_c)) when "00010000001", 
		    std_logic_vector(to_unsigned(878, n_bits_c)) when "00010000010", 
		    std_logic_vector(to_unsigned(880, n_bits_c)) when "00010000011", 
		    std_logic_vector(to_unsigned(881, n_bits_c)) when "00010000100", 
		    std_logic_vector(to_unsigned(883, n_bits_c)) when "00010000101", 
		    std_logic_vector(to_unsigned(885, n_bits_c)) when "00010000110", 
		    std_logic_vector(to_unsigned(886, n_bits_c)) when "00010000111", 
		    std_logic_vector(to_unsigned(888, n_bits_c)) when "00010001000", 
		    std_logic_vector(to_unsigned(889, n_bits_c)) when "00010001001", 
		    std_logic_vector(to_unsigned(891, n_bits_c)) when "00010001010", 
		    std_logic_vector(to_unsigned(892, n_bits_c)) when "00010001011", 
		    std_logic_vector(to_unsigned(894, n_bits_c)) when "00010001100", 
		    std_logic_vector(to_unsigned(895, n_bits_c)) when "00010001101", 
		    std_logic_vector(to_unsigned(897, n_bits_c)) when "00010001110", 
		    std_logic_vector(to_unsigned(898, n_bits_c)) when "00010001111", 
		    std_logic_vector(to_unsigned(900, n_bits_c)) when "00010010000", 
		    std_logic_vector(to_unsigned(901, n_bits_c)) when "00010010001", 
		    std_logic_vector(to_unsigned(903, n_bits_c)) when "00010010010", 
		    std_logic_vector(to_unsigned(904, n_bits_c)) when "00010010011", 
		    std_logic_vector(to_unsigned(906, n_bits_c)) when "00010010100", 
		    std_logic_vector(to_unsigned(907, n_bits_c)) when "00010010101", 
		    std_logic_vector(to_unsigned(909, n_bits_c)) when "00010010110", 
		    std_logic_vector(to_unsigned(910, n_bits_c)) when "00010010111", 
		    std_logic_vector(to_unsigned(912, n_bits_c)) when "00010011000", 
		    std_logic_vector(to_unsigned(913, n_bits_c)) when "00010011001", 
		    std_logic_vector(to_unsigned(915, n_bits_c)) when "00010011010", 
		    std_logic_vector(to_unsigned(916, n_bits_c)) when "00010011011", 
		    std_logic_vector(to_unsigned(918, n_bits_c)) when "00010011100", 
		    std_logic_vector(to_unsigned(919, n_bits_c)) when "00010011101", 
		    std_logic_vector(to_unsigned(921, n_bits_c)) when "00010011110", 
		    std_logic_vector(to_unsigned(922, n_bits_c)) when "00010011111", 
		    std_logic_vector(to_unsigned(924, n_bits_c)) when "00010100000", 
		    std_logic_vector(to_unsigned(925, n_bits_c)) when "00010100001", 
		    std_logic_vector(to_unsigned(926, n_bits_c)) when "00010100010", 
		    std_logic_vector(to_unsigned(928, n_bits_c)) when "00010100011", 
		    std_logic_vector(to_unsigned(929, n_bits_c)) when "00010100100", 
		    std_logic_vector(to_unsigned(931, n_bits_c)) when "00010100101", 
		    std_logic_vector(to_unsigned(932, n_bits_c)) when "00010100110", 
		    std_logic_vector(to_unsigned(934, n_bits_c)) when "00010100111", 
		    std_logic_vector(to_unsigned(935, n_bits_c)) when "00010101000", 
		    std_logic_vector(to_unsigned(937, n_bits_c)) when "00010101001", 
		    std_logic_vector(to_unsigned(938, n_bits_c)) when "00010101010", 
		    std_logic_vector(to_unsigned(940, n_bits_c)) when "00010101011", 
		    std_logic_vector(to_unsigned(941, n_bits_c)) when "00010101100", 
		    std_logic_vector(to_unsigned(942, n_bits_c)) when "00010101101", 
		    std_logic_vector(to_unsigned(944, n_bits_c)) when "00010101110", 
		    std_logic_vector(to_unsigned(945, n_bits_c)) when "00010101111", 
		    std_logic_vector(to_unsigned(947, n_bits_c)) when "00010110000", 
		    std_logic_vector(to_unsigned(948, n_bits_c)) when "00010110001", 
		    std_logic_vector(to_unsigned(950, n_bits_c)) when "00010110010", 
		    std_logic_vector(to_unsigned(951, n_bits_c)) when "00010110011", 
		    std_logic_vector(to_unsigned(952, n_bits_c)) when "00010110100", 
		    std_logic_vector(to_unsigned(954, n_bits_c)) when "00010110101", 
		    std_logic_vector(to_unsigned(955, n_bits_c)) when "00010110110", 
		    std_logic_vector(to_unsigned(957, n_bits_c)) when "00010110111", 
		    std_logic_vector(to_unsigned(958, n_bits_c)) when "00010111000", 
		    std_logic_vector(to_unsigned(959, n_bits_c)) when "00010111001", 
		    std_logic_vector(to_unsigned(961, n_bits_c)) when "00010111010", 
		    std_logic_vector(to_unsigned(962, n_bits_c)) when "00010111011", 
		    std_logic_vector(to_unsigned(964, n_bits_c)) when "00010111100", 
		    std_logic_vector(to_unsigned(965, n_bits_c)) when "00010111101", 
		    std_logic_vector(to_unsigned(966, n_bits_c)) when "00010111110", 
		    std_logic_vector(to_unsigned(968, n_bits_c)) when "00010111111", 
		    std_logic_vector(to_unsigned(969, n_bits_c)) when "00011000000", 
		    std_logic_vector(to_unsigned(971, n_bits_c)) when "00011000001", 
		    std_logic_vector(to_unsigned(972, n_bits_c)) when "00011000010", 
		    std_logic_vector(to_unsigned(973, n_bits_c)) when "00011000011", 
		    std_logic_vector(to_unsigned(975, n_bits_c)) when "00011000100", 
		    std_logic_vector(to_unsigned(976, n_bits_c)) when "00011000101", 
		    std_logic_vector(to_unsigned(978, n_bits_c)) when "00011000110", 
		    std_logic_vector(to_unsigned(979, n_bits_c)) when "00011000111", 
		    std_logic_vector(to_unsigned(980, n_bits_c)) when "00011001000", 
		    std_logic_vector(to_unsigned(982, n_bits_c)) when "00011001001", 
		    std_logic_vector(to_unsigned(983, n_bits_c)) when "00011001010", 
		    std_logic_vector(to_unsigned(984, n_bits_c)) when "00011001011", 
		    std_logic_vector(to_unsigned(986, n_bits_c)) when "00011001100", 
		    std_logic_vector(to_unsigned(987, n_bits_c)) when "00011001101", 
		    std_logic_vector(to_unsigned(988, n_bits_c)) when "00011001110", 
		    std_logic_vector(to_unsigned(990, n_bits_c)) when "00011001111", 
		    std_logic_vector(to_unsigned(991, n_bits_c)) when "00011010000", 
		    std_logic_vector(to_unsigned(992, n_bits_c)) when "00011010001", 
		    std_logic_vector(to_unsigned(994, n_bits_c)) when "00011010010", 
		    std_logic_vector(to_unsigned(995, n_bits_c)) when "00011010011", 
		    std_logic_vector(to_unsigned(996, n_bits_c)) when "00011010100", 
		    std_logic_vector(to_unsigned(998, n_bits_c)) when "00011010101", 
		    std_logic_vector(to_unsigned(999, n_bits_c)) when "00011010110", 
		    std_logic_vector(to_unsigned(1000, n_bits_c)) when "00011010111", 
		    std_logic_vector(to_unsigned(1002, n_bits_c)) when "00011011000", 
		    std_logic_vector(to_unsigned(1003, n_bits_c)) when "00011011001", 
		    std_logic_vector(to_unsigned(1004, n_bits_c)) when "00011011010", 
		    std_logic_vector(to_unsigned(1006, n_bits_c)) when "00011011011", 
		    std_logic_vector(to_unsigned(1007, n_bits_c)) when "00011011100", 
		    std_logic_vector(to_unsigned(1008, n_bits_c)) when "00011011101", 
		    std_logic_vector(to_unsigned(1009, n_bits_c)) when "00011011110", 
		    std_logic_vector(to_unsigned(1011, n_bits_c)) when "00011011111", 
		    std_logic_vector(to_unsigned(1012, n_bits_c)) when "00011100000", 
		    std_logic_vector(to_unsigned(1013, n_bits_c)) when "00011100001", 
		    std_logic_vector(to_unsigned(1015, n_bits_c)) when "00011100010", 
		    std_logic_vector(to_unsigned(1016, n_bits_c)) when "00011100011", 
		    std_logic_vector(to_unsigned(1017, n_bits_c)) when "00011100100", 
		    std_logic_vector(to_unsigned(1018, n_bits_c)) when "00011100101", 
		    std_logic_vector(to_unsigned(1020, n_bits_c)) when "00011100110", 
		    std_logic_vector(to_unsigned(1021, n_bits_c)) when "00011100111", 
		    std_logic_vector(to_unsigned(1022, n_bits_c)) when "00011101000", 
		    std_logic_vector(to_unsigned(1024, n_bits_c)) when "00011101001", 
		    std_logic_vector(to_unsigned(1025, n_bits_c)) when "00011101010", 
		    std_logic_vector(to_unsigned(1026, n_bits_c)) when "00011101011", 
		    std_logic_vector(to_unsigned(1027, n_bits_c)) when "00011101100", 
		    std_logic_vector(to_unsigned(1029, n_bits_c)) when "00011101101", 
		    std_logic_vector(to_unsigned(1030, n_bits_c)) when "00011101110", 
		    std_logic_vector(to_unsigned(1031, n_bits_c)) when "00011101111", 
		    std_logic_vector(to_unsigned(1032, n_bits_c)) when "00011110000", 
		    std_logic_vector(to_unsigned(1033, n_bits_c)) when "00011110001", 
		    std_logic_vector(to_unsigned(1035, n_bits_c)) when "00011110010", 
		    std_logic_vector(to_unsigned(1036, n_bits_c)) when "00011110011", 
		    std_logic_vector(to_unsigned(1037, n_bits_c)) when "00011110100", 
		    std_logic_vector(to_unsigned(1038, n_bits_c)) when "00011110101", 
		    std_logic_vector(to_unsigned(1040, n_bits_c)) when "00011110110", 
		    std_logic_vector(to_unsigned(1041, n_bits_c)) when "00011110111", 
		    std_logic_vector(to_unsigned(1042, n_bits_c)) when "00011111000", 
		    std_logic_vector(to_unsigned(1043, n_bits_c)) when "00011111001", 
		    std_logic_vector(to_unsigned(1044, n_bits_c)) when "00011111010", 
		    std_logic_vector(to_unsigned(1046, n_bits_c)) when "00011111011", 
		    std_logic_vector(to_unsigned(1047, n_bits_c)) when "00011111100", 
		    std_logic_vector(to_unsigned(1048, n_bits_c)) when "00011111101", 
		    std_logic_vector(to_unsigned(1049, n_bits_c)) when "00011111110", 
		    std_logic_vector(to_unsigned(1050, n_bits_c)) when "00011111111", 
		    std_logic_vector(to_unsigned(1052, n_bits_c)) when "00100000000", 
		    std_logic_vector(to_unsigned(1053, n_bits_c)) when "00100000001", 
		    std_logic_vector(to_unsigned(1054, n_bits_c)) when "00100000010", 
		    std_logic_vector(to_unsigned(1055, n_bits_c)) when "00100000011", 
		    std_logic_vector(to_unsigned(1056, n_bits_c)) when "00100000100", 
		    std_logic_vector(to_unsigned(1057, n_bits_c)) when "00100000101", 
		    std_logic_vector(to_unsigned(1059, n_bits_c)) when "00100000110", 
		    std_logic_vector(to_unsigned(1060, n_bits_c)) when "00100000111", 
		    std_logic_vector(to_unsigned(1061, n_bits_c)) when "00100001000", 
		    std_logic_vector(to_unsigned(1062, n_bits_c)) when "00100001001", 
		    std_logic_vector(to_unsigned(1063, n_bits_c)) when "00100001010", 
		    std_logic_vector(to_unsigned(1064, n_bits_c)) when "00100001011", 
		    std_logic_vector(to_unsigned(1065, n_bits_c)) when "00100001100", 
		    std_logic_vector(to_unsigned(1067, n_bits_c)) when "00100001101", 
		    std_logic_vector(to_unsigned(1068, n_bits_c)) when "00100001110", 
		    std_logic_vector(to_unsigned(1069, n_bits_c)) when "00100001111", 
		    std_logic_vector(to_unsigned(1070, n_bits_c)) when "00100010000", 
		    std_logic_vector(to_unsigned(1071, n_bits_c)) when "00100010001", 
		    std_logic_vector(to_unsigned(1072, n_bits_c)) when "00100010010", 
		    std_logic_vector(to_unsigned(1073, n_bits_c)) when "00100010011", 
		    std_logic_vector(to_unsigned(1074, n_bits_c)) when "00100010100", 
		    std_logic_vector(to_unsigned(1075, n_bits_c)) when "00100010101", 
		    std_logic_vector(to_unsigned(1077, n_bits_c)) when "00100010110", 
		    std_logic_vector(to_unsigned(1078, n_bits_c)) when "00100010111", 
		    std_logic_vector(to_unsigned(1079, n_bits_c)) when "00100011000", 
		    std_logic_vector(to_unsigned(1080, n_bits_c)) when "00100011001", 
		    std_logic_vector(to_unsigned(1081, n_bits_c)) when "00100011010", 
		    std_logic_vector(to_unsigned(1082, n_bits_c)) when "00100011011", 
		    std_logic_vector(to_unsigned(1083, n_bits_c)) when "00100011100", 
		    std_logic_vector(to_unsigned(1084, n_bits_c)) when "00100011101", 
		    std_logic_vector(to_unsigned(1085, n_bits_c)) when "00100011110", 
		    std_logic_vector(to_unsigned(1086, n_bits_c)) when "00100011111", 
		    std_logic_vector(to_unsigned(1087, n_bits_c)) when "00100100000", 
		    std_logic_vector(to_unsigned(1088, n_bits_c)) when "00100100001", 
		    std_logic_vector(to_unsigned(1089, n_bits_c)) when "00100100010", 
		    std_logic_vector(to_unsigned(1091, n_bits_c)) when "00100100011", 
		    std_logic_vector(to_unsigned(1092, n_bits_c)) when "00100100100", 
		    std_logic_vector(to_unsigned(1093, n_bits_c)) when "00100100101", 
		    std_logic_vector(to_unsigned(1094, n_bits_c)) when "00100100110", 
		    std_logic_vector(to_unsigned(1095, n_bits_c)) when "00100100111", 
		    std_logic_vector(to_unsigned(1096, n_bits_c)) when "00100101000", 
		    std_logic_vector(to_unsigned(1097, n_bits_c)) when "00100101001", 
		    std_logic_vector(to_unsigned(1098, n_bits_c)) when "00100101010", 
		    std_logic_vector(to_unsigned(1099, n_bits_c)) when "00100101011", 
		    std_logic_vector(to_unsigned(1100, n_bits_c)) when "00100101100", 
		    std_logic_vector(to_unsigned(1101, n_bits_c)) when "00100101101", 
		    std_logic_vector(to_unsigned(1102, n_bits_c)) when "00100101110", 
		    std_logic_vector(to_unsigned(1103, n_bits_c)) when "00100101111", 
		    std_logic_vector(to_unsigned(1104, n_bits_c)) when "00100110000", 
		    std_logic_vector(to_unsigned(1105, n_bits_c)) when "00100110001", 
		    std_logic_vector(to_unsigned(1106, n_bits_c)) when "00100110010", 
		    std_logic_vector(to_unsigned(1107, n_bits_c)) when "00100110011", 
		    std_logic_vector(to_unsigned(1108, n_bits_c)) when "00100110100", 
		    std_logic_vector(to_unsigned(1109, n_bits_c)) when "00100110101", 
		    std_logic_vector(to_unsigned(1110, n_bits_c)) when "00100110110", 
		    std_logic_vector(to_unsigned(1111, n_bits_c)) when "00100110111", 
		    std_logic_vector(to_unsigned(1112, n_bits_c)) when "00100111000", 
		    std_logic_vector(to_unsigned(1113, n_bits_c)) when "00100111001", 
		    std_logic_vector(to_unsigned(1113, n_bits_c)) when "00100111010", 
		    std_logic_vector(to_unsigned(1114, n_bits_c)) when "00100111011", 
		    std_logic_vector(to_unsigned(1115, n_bits_c)) when "00100111100", 
		    std_logic_vector(to_unsigned(1116, n_bits_c)) when "00100111101", 
		    std_logic_vector(to_unsigned(1117, n_bits_c)) when "00100111110", 
		    std_logic_vector(to_unsigned(1118, n_bits_c)) when "00100111111", 
		    std_logic_vector(to_unsigned(1119, n_bits_c)) when "00101000000", 
		    std_logic_vector(to_unsigned(1120, n_bits_c)) when "00101000001", 
		    std_logic_vector(to_unsigned(1121, n_bits_c)) when "00101000010", 
		    std_logic_vector(to_unsigned(1122, n_bits_c)) when "00101000011", 
		    std_logic_vector(to_unsigned(1123, n_bits_c)) when "00101000100", 
		    std_logic_vector(to_unsigned(1124, n_bits_c)) when "00101000101", 
		    std_logic_vector(to_unsigned(1125, n_bits_c)) when "00101000110", 
		    std_logic_vector(to_unsigned(1125, n_bits_c)) when "00101000111", 
		    std_logic_vector(to_unsigned(1126, n_bits_c)) when "00101001000", 
		    std_logic_vector(to_unsigned(1127, n_bits_c)) when "00101001001", 
		    std_logic_vector(to_unsigned(1128, n_bits_c)) when "00101001010", 
		    std_logic_vector(to_unsigned(1129, n_bits_c)) when "00101001011", 
		    std_logic_vector(to_unsigned(1130, n_bits_c)) when "00101001100", 
		    std_logic_vector(to_unsigned(1131, n_bits_c)) when "00101001101", 
		    std_logic_vector(to_unsigned(1132, n_bits_c)) when "00101001110", 
		    std_logic_vector(to_unsigned(1133, n_bits_c)) when "00101001111", 
		    std_logic_vector(to_unsigned(1133, n_bits_c)) when "00101010000", 
		    std_logic_vector(to_unsigned(1134, n_bits_c)) when "00101010001", 
		    std_logic_vector(to_unsigned(1135, n_bits_c)) when "00101010010", 
		    std_logic_vector(to_unsigned(1136, n_bits_c)) when "00101010011", 
		    std_logic_vector(to_unsigned(1137, n_bits_c)) when "00101010100", 
		    std_logic_vector(to_unsigned(1138, n_bits_c)) when "00101010101", 
		    std_logic_vector(to_unsigned(1138, n_bits_c)) when "00101010110", 
		    std_logic_vector(to_unsigned(1139, n_bits_c)) when "00101010111", 
		    std_logic_vector(to_unsigned(1140, n_bits_c)) when "00101011000", 
		    std_logic_vector(to_unsigned(1141, n_bits_c)) when "00101011001", 
		    std_logic_vector(to_unsigned(1142, n_bits_c)) when "00101011010", 
		    std_logic_vector(to_unsigned(1143, n_bits_c)) when "00101011011", 
		    std_logic_vector(to_unsigned(1143, n_bits_c)) when "00101011100", 
		    std_logic_vector(to_unsigned(1144, n_bits_c)) when "00101011101", 
		    std_logic_vector(to_unsigned(1145, n_bits_c)) when "00101011110", 
		    std_logic_vector(to_unsigned(1146, n_bits_c)) when "00101011111", 
		    std_logic_vector(to_unsigned(1147, n_bits_c)) when "00101100000", 
		    std_logic_vector(to_unsigned(1147, n_bits_c)) when "00101100001", 
		    std_logic_vector(to_unsigned(1148, n_bits_c)) when "00101100010", 
		    std_logic_vector(to_unsigned(1149, n_bits_c)) when "00101100011", 
		    std_logic_vector(to_unsigned(1150, n_bits_c)) when "00101100100", 
		    std_logic_vector(to_unsigned(1150, n_bits_c)) when "00101100101", 
		    std_logic_vector(to_unsigned(1151, n_bits_c)) when "00101100110", 
		    std_logic_vector(to_unsigned(1152, n_bits_c)) when "00101100111", 
		    std_logic_vector(to_unsigned(1153, n_bits_c)) when "00101101000", 
		    std_logic_vector(to_unsigned(1153, n_bits_c)) when "00101101001", 
		    std_logic_vector(to_unsigned(1154, n_bits_c)) when "00101101010", 
		    std_logic_vector(to_unsigned(1155, n_bits_c)) when "00101101011", 
		    std_logic_vector(to_unsigned(1156, n_bits_c)) when "00101101100", 
		    std_logic_vector(to_unsigned(1156, n_bits_c)) when "00101101101", 
		    std_logic_vector(to_unsigned(1157, n_bits_c)) when "00101101110", 
		    std_logic_vector(to_unsigned(1158, n_bits_c)) when "00101101111", 
		    std_logic_vector(to_unsigned(1158, n_bits_c)) when "00101110000", 
		    std_logic_vector(to_unsigned(1159, n_bits_c)) when "00101110001", 
		    std_logic_vector(to_unsigned(1160, n_bits_c)) when "00101110010", 
		    std_logic_vector(to_unsigned(1161, n_bits_c)) when "00101110011", 
		    std_logic_vector(to_unsigned(1161, n_bits_c)) when "00101110100", 
		    std_logic_vector(to_unsigned(1162, n_bits_c)) when "00101110101", 
		    std_logic_vector(to_unsigned(1163, n_bits_c)) when "00101110110", 
		    std_logic_vector(to_unsigned(1163, n_bits_c)) when "00101110111", 
		    std_logic_vector(to_unsigned(1164, n_bits_c)) when "00101111000", 
		    std_logic_vector(to_unsigned(1165, n_bits_c)) when "00101111001", 
		    std_logic_vector(to_unsigned(1165, n_bits_c)) when "00101111010", 
		    std_logic_vector(to_unsigned(1166, n_bits_c)) when "00101111011", 
		    std_logic_vector(to_unsigned(1167, n_bits_c)) when "00101111100", 
		    std_logic_vector(to_unsigned(1167, n_bits_c)) when "00101111101", 
		    std_logic_vector(to_unsigned(1168, n_bits_c)) when "00101111110", 
		    std_logic_vector(to_unsigned(1169, n_bits_c)) when "00101111111", 
		    std_logic_vector(to_unsigned(1169, n_bits_c)) when "00110000000", 
		    std_logic_vector(to_unsigned(1170, n_bits_c)) when "00110000001", 
		    std_logic_vector(to_unsigned(1171, n_bits_c)) when "00110000010", 
		    std_logic_vector(to_unsigned(1171, n_bits_c)) when "00110000011", 
		    std_logic_vector(to_unsigned(1172, n_bits_c)) when "00110000100", 
		    std_logic_vector(to_unsigned(1172, n_bits_c)) when "00110000101", 
		    std_logic_vector(to_unsigned(1173, n_bits_c)) when "00110000110", 
		    std_logic_vector(to_unsigned(1174, n_bits_c)) when "00110000111", 
		    std_logic_vector(to_unsigned(1174, n_bits_c)) when "00110001000", 
		    std_logic_vector(to_unsigned(1175, n_bits_c)) when "00110001001", 
		    std_logic_vector(to_unsigned(1175, n_bits_c)) when "00110001010", 
		    std_logic_vector(to_unsigned(1176, n_bits_c)) when "00110001011", 
		    std_logic_vector(to_unsigned(1177, n_bits_c)) when "00110001100", 
		    std_logic_vector(to_unsigned(1177, n_bits_c)) when "00110001101", 
		    std_logic_vector(to_unsigned(1178, n_bits_c)) when "00110001110", 
		    std_logic_vector(to_unsigned(1178, n_bits_c)) when "00110001111", 
		    std_logic_vector(to_unsigned(1179, n_bits_c)) when "00110010000", 
		    std_logic_vector(to_unsigned(1179, n_bits_c)) when "00110010001", 
		    std_logic_vector(to_unsigned(1180, n_bits_c)) when "00110010010", 
		    std_logic_vector(to_unsigned(1181, n_bits_c)) when "00110010011", 
		    std_logic_vector(to_unsigned(1181, n_bits_c)) when "00110010100", 
		    std_logic_vector(to_unsigned(1182, n_bits_c)) when "00110010101", 
		    std_logic_vector(to_unsigned(1182, n_bits_c)) when "00110010110", 
		    std_logic_vector(to_unsigned(1183, n_bits_c)) when "00110010111", 
		    std_logic_vector(to_unsigned(1183, n_bits_c)) when "00110011000", 
		    std_logic_vector(to_unsigned(1184, n_bits_c)) when "00110011001", 
		    std_logic_vector(to_unsigned(1184, n_bits_c)) when "00110011010", 
		    std_logic_vector(to_unsigned(1185, n_bits_c)) when "00110011011", 
		    std_logic_vector(to_unsigned(1185, n_bits_c)) when "00110011100", 
		    std_logic_vector(to_unsigned(1186, n_bits_c)) when "00110011101", 
		    std_logic_vector(to_unsigned(1186, n_bits_c)) when "00110011110", 
		    std_logic_vector(to_unsigned(1187, n_bits_c)) when "00110011111", 
		    std_logic_vector(to_unsigned(1187, n_bits_c)) when "00110100000", 
		    std_logic_vector(to_unsigned(1188, n_bits_c)) when "00110100001", 
		    std_logic_vector(to_unsigned(1188, n_bits_c)) when "00110100010", 
		    std_logic_vector(to_unsigned(1189, n_bits_c)) when "00110100011", 
		    std_logic_vector(to_unsigned(1189, n_bits_c)) when "00110100100", 
		    std_logic_vector(to_unsigned(1190, n_bits_c)) when "00110100101", 
		    std_logic_vector(to_unsigned(1190, n_bits_c)) when "00110100110", 
		    std_logic_vector(to_unsigned(1191, n_bits_c)) when "00110100111", 
		    std_logic_vector(to_unsigned(1191, n_bits_c)) when "00110101000", 
		    std_logic_vector(to_unsigned(1191, n_bits_c)) when "00110101001", 
		    std_logic_vector(to_unsigned(1192, n_bits_c)) when "00110101010", 
		    std_logic_vector(to_unsigned(1192, n_bits_c)) when "00110101011", 
		    std_logic_vector(to_unsigned(1193, n_bits_c)) when "00110101100", 
		    std_logic_vector(to_unsigned(1193, n_bits_c)) when "00110101101", 
		    std_logic_vector(to_unsigned(1194, n_bits_c)) when "00110101110", 
		    std_logic_vector(to_unsigned(1194, n_bits_c)) when "00110101111", 
		    std_logic_vector(to_unsigned(1194, n_bits_c)) when "00110110000", 
		    std_logic_vector(to_unsigned(1195, n_bits_c)) when "00110110001", 
		    std_logic_vector(to_unsigned(1195, n_bits_c)) when "00110110010", 
		    std_logic_vector(to_unsigned(1196, n_bits_c)) when "00110110011", 
		    std_logic_vector(to_unsigned(1196, n_bits_c)) when "00110110100", 
		    std_logic_vector(to_unsigned(1196, n_bits_c)) when "00110110101", 
		    std_logic_vector(to_unsigned(1197, n_bits_c)) when "00110110110", 
		    std_logic_vector(to_unsigned(1197, n_bits_c)) when "00110110111", 
		    std_logic_vector(to_unsigned(1197, n_bits_c)) when "00110111000", 
		    std_logic_vector(to_unsigned(1198, n_bits_c)) when "00110111001", 
		    std_logic_vector(to_unsigned(1198, n_bits_c)) when "00110111010", 
		    std_logic_vector(to_unsigned(1199, n_bits_c)) when "00110111011", 
		    std_logic_vector(to_unsigned(1199, n_bits_c)) when "00110111100", 
		    std_logic_vector(to_unsigned(1199, n_bits_c)) when "00110111101", 
		    std_logic_vector(to_unsigned(1200, n_bits_c)) when "00110111110", 
		    std_logic_vector(to_unsigned(1200, n_bits_c)) when "00110111111", 
		    std_logic_vector(to_unsigned(1200, n_bits_c)) when "00111000000", 
		    std_logic_vector(to_unsigned(1201, n_bits_c)) when "00111000001", 
		    std_logic_vector(to_unsigned(1201, n_bits_c)) when "00111000010", 
		    std_logic_vector(to_unsigned(1201, n_bits_c)) when "00111000011", 
		    std_logic_vector(to_unsigned(1201, n_bits_c)) when "00111000100", 
		    std_logic_vector(to_unsigned(1202, n_bits_c)) when "00111000101", 
		    std_logic_vector(to_unsigned(1202, n_bits_c)) when "00111000110", 
		    std_logic_vector(to_unsigned(1202, n_bits_c)) when "00111000111", 
		    std_logic_vector(to_unsigned(1203, n_bits_c)) when "00111001000", 
		    std_logic_vector(to_unsigned(1203, n_bits_c)) when "00111001001", 
		    std_logic_vector(to_unsigned(1203, n_bits_c)) when "00111001010", 
		    std_logic_vector(to_unsigned(1203, n_bits_c)) when "00111001011", 
		    std_logic_vector(to_unsigned(1204, n_bits_c)) when "00111001100", 
		    std_logic_vector(to_unsigned(1204, n_bits_c)) when "00111001101", 
		    std_logic_vector(to_unsigned(1204, n_bits_c)) when "00111001110", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "00111001111", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "00111010000", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "00111010001", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "00111010010", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "00111010011", 
		    std_logic_vector(to_unsigned(1206, n_bits_c)) when "00111010100", 
		    std_logic_vector(to_unsigned(1206, n_bits_c)) when "00111010101", 
		    std_logic_vector(to_unsigned(1206, n_bits_c)) when "00111010110", 
		    std_logic_vector(to_unsigned(1206, n_bits_c)) when "00111010111", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "00111011000", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "00111011001", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "00111011010", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "00111011011", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "00111011100", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "00111011101", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "00111011110", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "00111011111", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "00111100000", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "00111100001", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "00111100010", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "00111100011", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "00111100100", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "00111100101", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "00111100110", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "00111100111", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "00111101000", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "00111101001", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "00111101010", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111101011", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111101100", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111101101", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111101110", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111101111", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111110000", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111110001", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111110010", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111110011", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111110100", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111110101", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111110110", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111110111", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "00111111000", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "00111111001", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "00111111010", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "00111111011", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "00111111100", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "00111111101", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "00111111110", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "00111111111", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "01000000000", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "01000000001", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "01000000010", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "01000000011", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "01000000100", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "01000000101", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "01000000110", 
		    std_logic_vector(to_unsigned(1211, n_bits_c)) when "01000000111", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000001000", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000001001", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000001010", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000001011", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000001100", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000001101", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000001110", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000001111", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000010000", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000010001", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000010010", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000010011", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000010100", 
		    std_logic_vector(to_unsigned(1210, n_bits_c)) when "01000010101", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "01000010110", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "01000010111", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "01000011000", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "01000011001", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "01000011010", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "01000011011", 
		    std_logic_vector(to_unsigned(1209, n_bits_c)) when "01000011100", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "01000011101", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "01000011110", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "01000011111", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "01000100000", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "01000100001", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "01000100010", 
		    std_logic_vector(to_unsigned(1208, n_bits_c)) when "01000100011", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "01000100100", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "01000100101", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "01000100110", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "01000100111", 
		    std_logic_vector(to_unsigned(1207, n_bits_c)) when "01000101000", 
		    std_logic_vector(to_unsigned(1206, n_bits_c)) when "01000101001", 
		    std_logic_vector(to_unsigned(1206, n_bits_c)) when "01000101010", 
		    std_logic_vector(to_unsigned(1206, n_bits_c)) when "01000101011", 
		    std_logic_vector(to_unsigned(1206, n_bits_c)) when "01000101100", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "01000101101", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "01000101110", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "01000101111", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "01000110000", 
		    std_logic_vector(to_unsigned(1205, n_bits_c)) when "01000110001", 
		    std_logic_vector(to_unsigned(1204, n_bits_c)) when "01000110010", 
		    std_logic_vector(to_unsigned(1204, n_bits_c)) when "01000110011", 
		    std_logic_vector(to_unsigned(1204, n_bits_c)) when "01000110100", 
		    std_logic_vector(to_unsigned(1203, n_bits_c)) when "01000110101", 
		    std_logic_vector(to_unsigned(1203, n_bits_c)) when "01000110110", 
		    std_logic_vector(to_unsigned(1203, n_bits_c)) when "01000110111", 
		    std_logic_vector(to_unsigned(1203, n_bits_c)) when "01000111000", 
		    std_logic_vector(to_unsigned(1202, n_bits_c)) when "01000111001", 
		    std_logic_vector(to_unsigned(1202, n_bits_c)) when "01000111010", 
		    std_logic_vector(to_unsigned(1202, n_bits_c)) when "01000111011", 
		    std_logic_vector(to_unsigned(1201, n_bits_c)) when "01000111100", 
		    std_logic_vector(to_unsigned(1201, n_bits_c)) when "01000111101", 
		    std_logic_vector(to_unsigned(1201, n_bits_c)) when "01000111110", 
		    std_logic_vector(to_unsigned(1201, n_bits_c)) when "01000111111", 
		    std_logic_vector(to_unsigned(1200, n_bits_c)) when "01001000000", 
		    std_logic_vector(to_unsigned(1200, n_bits_c)) when "01001000001", 
		    std_logic_vector(to_unsigned(1200, n_bits_c)) when "01001000010", 
		    std_logic_vector(to_unsigned(1199, n_bits_c)) when "01001000011", 
		    std_logic_vector(to_unsigned(1199, n_bits_c)) when "01001000100", 
		    std_logic_vector(to_unsigned(1199, n_bits_c)) when "01001000101", 
		    std_logic_vector(to_unsigned(1198, n_bits_c)) when "01001000110", 
		    std_logic_vector(to_unsigned(1198, n_bits_c)) when "01001000111", 
		    std_logic_vector(to_unsigned(1197, n_bits_c)) when "01001001000", 
		    std_logic_vector(to_unsigned(1197, n_bits_c)) when "01001001001", 
		    std_logic_vector(to_unsigned(1197, n_bits_c)) when "01001001010", 
		    std_logic_vector(to_unsigned(1196, n_bits_c)) when "01001001011", 
		    std_logic_vector(to_unsigned(1196, n_bits_c)) when "01001001100", 
		    std_logic_vector(to_unsigned(1196, n_bits_c)) when "01001001101", 
		    std_logic_vector(to_unsigned(1195, n_bits_c)) when "01001001110", 
		    std_logic_vector(to_unsigned(1195, n_bits_c)) when "01001001111", 
		    std_logic_vector(to_unsigned(1194, n_bits_c)) when "01001010000", 
		    std_logic_vector(to_unsigned(1194, n_bits_c)) when "01001010001", 
		    std_logic_vector(to_unsigned(1194, n_bits_c)) when "01001010010", 
		    std_logic_vector(to_unsigned(1193, n_bits_c)) when "01001010011", 
		    std_logic_vector(to_unsigned(1193, n_bits_c)) when "01001010100", 
		    std_logic_vector(to_unsigned(1192, n_bits_c)) when "01001010101", 
		    std_logic_vector(to_unsigned(1192, n_bits_c)) when "01001010110", 
		    std_logic_vector(to_unsigned(1191, n_bits_c)) when "01001010111", 
		    std_logic_vector(to_unsigned(1191, n_bits_c)) when "01001011000", 
		    std_logic_vector(to_unsigned(1191, n_bits_c)) when "01001011001", 
		    std_logic_vector(to_unsigned(1190, n_bits_c)) when "01001011010", 
		    std_logic_vector(to_unsigned(1190, n_bits_c)) when "01001011011", 
		    std_logic_vector(to_unsigned(1189, n_bits_c)) when "01001011100", 
		    std_logic_vector(to_unsigned(1189, n_bits_c)) when "01001011101", 
		    std_logic_vector(to_unsigned(1188, n_bits_c)) when "01001011110", 
		    std_logic_vector(to_unsigned(1188, n_bits_c)) when "01001011111", 
		    std_logic_vector(to_unsigned(1187, n_bits_c)) when "01001100000", 
		    std_logic_vector(to_unsigned(1187, n_bits_c)) when "01001100001", 
		    std_logic_vector(to_unsigned(1186, n_bits_c)) when "01001100010", 
		    std_logic_vector(to_unsigned(1186, n_bits_c)) when "01001100011", 
		    std_logic_vector(to_unsigned(1185, n_bits_c)) when "01001100100", 
		    std_logic_vector(to_unsigned(1185, n_bits_c)) when "01001100101", 
		    std_logic_vector(to_unsigned(1184, n_bits_c)) when "01001100110", 
		    std_logic_vector(to_unsigned(1184, n_bits_c)) when "01001100111", 
		    std_logic_vector(to_unsigned(1183, n_bits_c)) when "01001101000", 
		    std_logic_vector(to_unsigned(1183, n_bits_c)) when "01001101001", 
		    std_logic_vector(to_unsigned(1182, n_bits_c)) when "01001101010", 
		    std_logic_vector(to_unsigned(1182, n_bits_c)) when "01001101011", 
		    std_logic_vector(to_unsigned(1181, n_bits_c)) when "01001101100", 
		    std_logic_vector(to_unsigned(1181, n_bits_c)) when "01001101101", 
		    std_logic_vector(to_unsigned(1180, n_bits_c)) when "01001101110", 
		    std_logic_vector(to_unsigned(1179, n_bits_c)) when "01001101111", 
		    std_logic_vector(to_unsigned(1179, n_bits_c)) when "01001110000", 
		    std_logic_vector(to_unsigned(1178, n_bits_c)) when "01001110001", 
		    std_logic_vector(to_unsigned(1178, n_bits_c)) when "01001110010", 
		    std_logic_vector(to_unsigned(1177, n_bits_c)) when "01001110011", 
		    std_logic_vector(to_unsigned(1177, n_bits_c)) when "01001110100", 
		    std_logic_vector(to_unsigned(1176, n_bits_c)) when "01001110101", 
		    std_logic_vector(to_unsigned(1175, n_bits_c)) when "01001110110", 
		    std_logic_vector(to_unsigned(1175, n_bits_c)) when "01001110111", 
		    std_logic_vector(to_unsigned(1174, n_bits_c)) when "01001111000", 
		    std_logic_vector(to_unsigned(1174, n_bits_c)) when "01001111001", 
		    std_logic_vector(to_unsigned(1173, n_bits_c)) when "01001111010", 
		    std_logic_vector(to_unsigned(1172, n_bits_c)) when "01001111011", 
		    std_logic_vector(to_unsigned(1172, n_bits_c)) when "01001111100", 
		    std_logic_vector(to_unsigned(1171, n_bits_c)) when "01001111101", 
		    std_logic_vector(to_unsigned(1171, n_bits_c)) when "01001111110", 
		    std_logic_vector(to_unsigned(1170, n_bits_c)) when "01001111111", 
		    std_logic_vector(to_unsigned(1169, n_bits_c)) when "01010000000", 
		    std_logic_vector(to_unsigned(1169, n_bits_c)) when "01010000001", 
		    std_logic_vector(to_unsigned(1168, n_bits_c)) when "01010000010", 
		    std_logic_vector(to_unsigned(1167, n_bits_c)) when "01010000011", 
		    std_logic_vector(to_unsigned(1167, n_bits_c)) when "01010000100", 
		    std_logic_vector(to_unsigned(1166, n_bits_c)) when "01010000101", 
		    std_logic_vector(to_unsigned(1165, n_bits_c)) when "01010000110", 
		    std_logic_vector(to_unsigned(1165, n_bits_c)) when "01010000111", 
		    std_logic_vector(to_unsigned(1164, n_bits_c)) when "01010001000", 
		    std_logic_vector(to_unsigned(1163, n_bits_c)) when "01010001001", 
		    std_logic_vector(to_unsigned(1163, n_bits_c)) when "01010001010", 
		    std_logic_vector(to_unsigned(1162, n_bits_c)) when "01010001011", 
		    std_logic_vector(to_unsigned(1161, n_bits_c)) when "01010001100", 
		    std_logic_vector(to_unsigned(1161, n_bits_c)) when "01010001101", 
		    std_logic_vector(to_unsigned(1160, n_bits_c)) when "01010001110", 
		    std_logic_vector(to_unsigned(1159, n_bits_c)) when "01010001111", 
		    std_logic_vector(to_unsigned(1158, n_bits_c)) when "01010010000", 
		    std_logic_vector(to_unsigned(1158, n_bits_c)) when "01010010001", 
		    std_logic_vector(to_unsigned(1157, n_bits_c)) when "01010010010", 
		    std_logic_vector(to_unsigned(1156, n_bits_c)) when "01010010011", 
		    std_logic_vector(to_unsigned(1156, n_bits_c)) when "01010010100", 
		    std_logic_vector(to_unsigned(1155, n_bits_c)) when "01010010101", 
		    std_logic_vector(to_unsigned(1154, n_bits_c)) when "01010010110", 
		    std_logic_vector(to_unsigned(1153, n_bits_c)) when "01010010111", 
		    std_logic_vector(to_unsigned(1153, n_bits_c)) when "01010011000", 
		    std_logic_vector(to_unsigned(1152, n_bits_c)) when "01010011001", 
		    std_logic_vector(to_unsigned(1151, n_bits_c)) when "01010011010", 
		    std_logic_vector(to_unsigned(1150, n_bits_c)) when "01010011011", 
		    std_logic_vector(to_unsigned(1150, n_bits_c)) when "01010011100", 
		    std_logic_vector(to_unsigned(1149, n_bits_c)) when "01010011101", 
		    std_logic_vector(to_unsigned(1148, n_bits_c)) when "01010011110", 
		    std_logic_vector(to_unsigned(1147, n_bits_c)) when "01010011111", 
		    std_logic_vector(to_unsigned(1147, n_bits_c)) when "01010100000", 
		    std_logic_vector(to_unsigned(1146, n_bits_c)) when "01010100001", 
		    std_logic_vector(to_unsigned(1145, n_bits_c)) when "01010100010", 
		    std_logic_vector(to_unsigned(1144, n_bits_c)) when "01010100011", 
		    std_logic_vector(to_unsigned(1143, n_bits_c)) when "01010100100", 
		    std_logic_vector(to_unsigned(1143, n_bits_c)) when "01010100101", 
		    std_logic_vector(to_unsigned(1142, n_bits_c)) when "01010100110", 
		    std_logic_vector(to_unsigned(1141, n_bits_c)) when "01010100111", 
		    std_logic_vector(to_unsigned(1140, n_bits_c)) when "01010101000", 
		    std_logic_vector(to_unsigned(1139, n_bits_c)) when "01010101001", 
		    std_logic_vector(to_unsigned(1138, n_bits_c)) when "01010101010", 
		    std_logic_vector(to_unsigned(1138, n_bits_c)) when "01010101011", 
		    std_logic_vector(to_unsigned(1137, n_bits_c)) when "01010101100", 
		    std_logic_vector(to_unsigned(1136, n_bits_c)) when "01010101101", 
		    std_logic_vector(to_unsigned(1135, n_bits_c)) when "01010101110", 
		    std_logic_vector(to_unsigned(1134, n_bits_c)) when "01010101111", 
		    std_logic_vector(to_unsigned(1133, n_bits_c)) when "01010110000", 
		    std_logic_vector(to_unsigned(1133, n_bits_c)) when "01010110001", 
		    std_logic_vector(to_unsigned(1132, n_bits_c)) when "01010110010", 
		    std_logic_vector(to_unsigned(1131, n_bits_c)) when "01010110011", 
		    std_logic_vector(to_unsigned(1130, n_bits_c)) when "01010110100", 
		    std_logic_vector(to_unsigned(1129, n_bits_c)) when "01010110101", 
		    std_logic_vector(to_unsigned(1128, n_bits_c)) when "01010110110", 
		    std_logic_vector(to_unsigned(1127, n_bits_c)) when "01010110111", 
		    std_logic_vector(to_unsigned(1126, n_bits_c)) when "01010111000", 
		    std_logic_vector(to_unsigned(1125, n_bits_c)) when "01010111001", 
		    std_logic_vector(to_unsigned(1125, n_bits_c)) when "01010111010", 
		    std_logic_vector(to_unsigned(1124, n_bits_c)) when "01010111011", 
		    std_logic_vector(to_unsigned(1123, n_bits_c)) when "01010111100", 
		    std_logic_vector(to_unsigned(1122, n_bits_c)) when "01010111101", 
		    std_logic_vector(to_unsigned(1121, n_bits_c)) when "01010111110", 
		    std_logic_vector(to_unsigned(1120, n_bits_c)) when "01010111111", 
		    std_logic_vector(to_unsigned(1119, n_bits_c)) when "01011000000", 
		    std_logic_vector(to_unsigned(1118, n_bits_c)) when "01011000001", 
		    std_logic_vector(to_unsigned(1117, n_bits_c)) when "01011000010", 
		    std_logic_vector(to_unsigned(1116, n_bits_c)) when "01011000011", 
		    std_logic_vector(to_unsigned(1115, n_bits_c)) when "01011000100", 
		    std_logic_vector(to_unsigned(1114, n_bits_c)) when "01011000101", 
		    std_logic_vector(to_unsigned(1113, n_bits_c)) when "01011000110", 
		    std_logic_vector(to_unsigned(1113, n_bits_c)) when "01011000111", 
		    std_logic_vector(to_unsigned(1112, n_bits_c)) when "01011001000", 
		    std_logic_vector(to_unsigned(1111, n_bits_c)) when "01011001001", 
		    std_logic_vector(to_unsigned(1110, n_bits_c)) when "01011001010", 
		    std_logic_vector(to_unsigned(1109, n_bits_c)) when "01011001011", 
		    std_logic_vector(to_unsigned(1108, n_bits_c)) when "01011001100", 
		    std_logic_vector(to_unsigned(1107, n_bits_c)) when "01011001101", 
		    std_logic_vector(to_unsigned(1106, n_bits_c)) when "01011001110", 
		    std_logic_vector(to_unsigned(1105, n_bits_c)) when "01011001111", 
		    std_logic_vector(to_unsigned(1104, n_bits_c)) when "01011010000", 
		    std_logic_vector(to_unsigned(1103, n_bits_c)) when "01011010001", 
		    std_logic_vector(to_unsigned(1102, n_bits_c)) when "01011010010", 
		    std_logic_vector(to_unsigned(1101, n_bits_c)) when "01011010011", 
		    std_logic_vector(to_unsigned(1100, n_bits_c)) when "01011010100", 
		    std_logic_vector(to_unsigned(1099, n_bits_c)) when "01011010101", 
		    std_logic_vector(to_unsigned(1098, n_bits_c)) when "01011010110", 
		    std_logic_vector(to_unsigned(1097, n_bits_c)) when "01011010111", 
		    std_logic_vector(to_unsigned(1096, n_bits_c)) when "01011011000", 
		    std_logic_vector(to_unsigned(1095, n_bits_c)) when "01011011001", 
		    std_logic_vector(to_unsigned(1094, n_bits_c)) when "01011011010", 
		    std_logic_vector(to_unsigned(1093, n_bits_c)) when "01011011011", 
		    std_logic_vector(to_unsigned(1092, n_bits_c)) when "01011011100", 
		    std_logic_vector(to_unsigned(1091, n_bits_c)) when "01011011101", 
		    std_logic_vector(to_unsigned(1089, n_bits_c)) when "01011011110", 
		    std_logic_vector(to_unsigned(1088, n_bits_c)) when "01011011111", 
		    std_logic_vector(to_unsigned(1087, n_bits_c)) when "01011100000", 
		    std_logic_vector(to_unsigned(1086, n_bits_c)) when "01011100001", 
		    std_logic_vector(to_unsigned(1085, n_bits_c)) when "01011100010", 
		    std_logic_vector(to_unsigned(1084, n_bits_c)) when "01011100011", 
		    std_logic_vector(to_unsigned(1083, n_bits_c)) when "01011100100", 
		    std_logic_vector(to_unsigned(1082, n_bits_c)) when "01011100101", 
		    std_logic_vector(to_unsigned(1081, n_bits_c)) when "01011100110", 
		    std_logic_vector(to_unsigned(1080, n_bits_c)) when "01011100111", 
		    std_logic_vector(to_unsigned(1079, n_bits_c)) when "01011101000", 
		    std_logic_vector(to_unsigned(1078, n_bits_c)) when "01011101001", 
		    std_logic_vector(to_unsigned(1077, n_bits_c)) when "01011101010", 
		    std_logic_vector(to_unsigned(1075, n_bits_c)) when "01011101011", 
		    std_logic_vector(to_unsigned(1074, n_bits_c)) when "01011101100", 
		    std_logic_vector(to_unsigned(1073, n_bits_c)) when "01011101101", 
		    std_logic_vector(to_unsigned(1072, n_bits_c)) when "01011101110", 
		    std_logic_vector(to_unsigned(1071, n_bits_c)) when "01011101111", 
		    std_logic_vector(to_unsigned(1070, n_bits_c)) when "01011110000", 
		    std_logic_vector(to_unsigned(1069, n_bits_c)) when "01011110001", 
		    std_logic_vector(to_unsigned(1068, n_bits_c)) when "01011110010", 
		    std_logic_vector(to_unsigned(1067, n_bits_c)) when "01011110011", 
		    std_logic_vector(to_unsigned(1065, n_bits_c)) when "01011110100", 
		    std_logic_vector(to_unsigned(1064, n_bits_c)) when "01011110101", 
		    std_logic_vector(to_unsigned(1063, n_bits_c)) when "01011110110", 
		    std_logic_vector(to_unsigned(1062, n_bits_c)) when "01011110111", 
		    std_logic_vector(to_unsigned(1061, n_bits_c)) when "01011111000", 
		    std_logic_vector(to_unsigned(1060, n_bits_c)) when "01011111001", 
		    std_logic_vector(to_unsigned(1059, n_bits_c)) when "01011111010", 
		    std_logic_vector(to_unsigned(1057, n_bits_c)) when "01011111011", 
		    std_logic_vector(to_unsigned(1056, n_bits_c)) when "01011111100", 
		    std_logic_vector(to_unsigned(1055, n_bits_c)) when "01011111101", 
		    std_logic_vector(to_unsigned(1054, n_bits_c)) when "01011111110", 
		    std_logic_vector(to_unsigned(1053, n_bits_c)) when "01011111111", 
		    std_logic_vector(to_unsigned(1052, n_bits_c)) when "01100000000", 
		    std_logic_vector(to_unsigned(1050, n_bits_c)) when "01100000001", 
		    std_logic_vector(to_unsigned(1049, n_bits_c)) when "01100000010", 
		    std_logic_vector(to_unsigned(1048, n_bits_c)) when "01100000011", 
		    std_logic_vector(to_unsigned(1047, n_bits_c)) when "01100000100", 
		    std_logic_vector(to_unsigned(1046, n_bits_c)) when "01100000101", 
		    std_logic_vector(to_unsigned(1044, n_bits_c)) when "01100000110", 
		    std_logic_vector(to_unsigned(1043, n_bits_c)) when "01100000111", 
		    std_logic_vector(to_unsigned(1042, n_bits_c)) when "01100001000", 
		    std_logic_vector(to_unsigned(1041, n_bits_c)) when "01100001001", 
		    std_logic_vector(to_unsigned(1040, n_bits_c)) when "01100001010", 
		    std_logic_vector(to_unsigned(1038, n_bits_c)) when "01100001011", 
		    std_logic_vector(to_unsigned(1037, n_bits_c)) when "01100001100", 
		    std_logic_vector(to_unsigned(1036, n_bits_c)) when "01100001101", 
		    std_logic_vector(to_unsigned(1035, n_bits_c)) when "01100001110", 
		    std_logic_vector(to_unsigned(1033, n_bits_c)) when "01100001111", 
		    std_logic_vector(to_unsigned(1032, n_bits_c)) when "01100010000", 
		    std_logic_vector(to_unsigned(1031, n_bits_c)) when "01100010001", 
		    std_logic_vector(to_unsigned(1030, n_bits_c)) when "01100010010", 
		    std_logic_vector(to_unsigned(1029, n_bits_c)) when "01100010011", 
		    std_logic_vector(to_unsigned(1027, n_bits_c)) when "01100010100", 
		    std_logic_vector(to_unsigned(1026, n_bits_c)) when "01100010101", 
		    std_logic_vector(to_unsigned(1025, n_bits_c)) when "01100010110", 
		    std_logic_vector(to_unsigned(1024, n_bits_c)) when "01100010111", 
		    std_logic_vector(to_unsigned(1022, n_bits_c)) when "01100011000", 
		    std_logic_vector(to_unsigned(1021, n_bits_c)) when "01100011001", 
		    std_logic_vector(to_unsigned(1020, n_bits_c)) when "01100011010", 
		    std_logic_vector(to_unsigned(1018, n_bits_c)) when "01100011011", 
		    std_logic_vector(to_unsigned(1017, n_bits_c)) when "01100011100", 
		    std_logic_vector(to_unsigned(1016, n_bits_c)) when "01100011101", 
		    std_logic_vector(to_unsigned(1015, n_bits_c)) when "01100011110", 
		    std_logic_vector(to_unsigned(1013, n_bits_c)) when "01100011111", 
		    std_logic_vector(to_unsigned(1012, n_bits_c)) when "01100100000", 
		    std_logic_vector(to_unsigned(1011, n_bits_c)) when "01100100001", 
		    std_logic_vector(to_unsigned(1009, n_bits_c)) when "01100100010", 
		    std_logic_vector(to_unsigned(1008, n_bits_c)) when "01100100011", 
		    std_logic_vector(to_unsigned(1007, n_bits_c)) when "01100100100", 
		    std_logic_vector(to_unsigned(1006, n_bits_c)) when "01100100101", 
		    std_logic_vector(to_unsigned(1004, n_bits_c)) when "01100100110", 
		    std_logic_vector(to_unsigned(1003, n_bits_c)) when "01100100111", 
		    std_logic_vector(to_unsigned(1002, n_bits_c)) when "01100101000", 
		    std_logic_vector(to_unsigned(1000, n_bits_c)) when "01100101001", 
		    std_logic_vector(to_unsigned(999, n_bits_c)) when "01100101010", 
		    std_logic_vector(to_unsigned(998, n_bits_c)) when "01100101011", 
		    std_logic_vector(to_unsigned(996, n_bits_c)) when "01100101100", 
		    std_logic_vector(to_unsigned(995, n_bits_c)) when "01100101101", 
		    std_logic_vector(to_unsigned(994, n_bits_c)) when "01100101110", 
		    std_logic_vector(to_unsigned(992, n_bits_c)) when "01100101111", 
		    std_logic_vector(to_unsigned(991, n_bits_c)) when "01100110000", 
		    std_logic_vector(to_unsigned(990, n_bits_c)) when "01100110001", 
		    std_logic_vector(to_unsigned(988, n_bits_c)) when "01100110010", 
		    std_logic_vector(to_unsigned(987, n_bits_c)) when "01100110011", 
		    std_logic_vector(to_unsigned(986, n_bits_c)) when "01100110100", 
		    std_logic_vector(to_unsigned(984, n_bits_c)) when "01100110101", 
		    std_logic_vector(to_unsigned(983, n_bits_c)) when "01100110110", 
		    std_logic_vector(to_unsigned(982, n_bits_c)) when "01100110111", 
		    std_logic_vector(to_unsigned(980, n_bits_c)) when "01100111000", 
		    std_logic_vector(to_unsigned(979, n_bits_c)) when "01100111001", 
		    std_logic_vector(to_unsigned(978, n_bits_c)) when "01100111010", 
		    std_logic_vector(to_unsigned(976, n_bits_c)) when "01100111011", 
		    std_logic_vector(to_unsigned(975, n_bits_c)) when "01100111100", 
		    std_logic_vector(to_unsigned(973, n_bits_c)) when "01100111101", 
		    std_logic_vector(to_unsigned(972, n_bits_c)) when "01100111110", 
		    std_logic_vector(to_unsigned(971, n_bits_c)) when "01100111111", 
		    std_logic_vector(to_unsigned(969, n_bits_c)) when "01101000000", 
		    std_logic_vector(to_unsigned(968, n_bits_c)) when "01101000001", 
		    std_logic_vector(to_unsigned(966, n_bits_c)) when "01101000010", 
		    std_logic_vector(to_unsigned(965, n_bits_c)) when "01101000011", 
		    std_logic_vector(to_unsigned(964, n_bits_c)) when "01101000100", 
		    std_logic_vector(to_unsigned(962, n_bits_c)) when "01101000101", 
		    std_logic_vector(to_unsigned(961, n_bits_c)) when "01101000110", 
		    std_logic_vector(to_unsigned(959, n_bits_c)) when "01101000111", 
		    std_logic_vector(to_unsigned(958, n_bits_c)) when "01101001000", 
		    std_logic_vector(to_unsigned(957, n_bits_c)) when "01101001001", 
		    std_logic_vector(to_unsigned(955, n_bits_c)) when "01101001010", 
		    std_logic_vector(to_unsigned(954, n_bits_c)) when "01101001011", 
		    std_logic_vector(to_unsigned(952, n_bits_c)) when "01101001100", 
		    std_logic_vector(to_unsigned(951, n_bits_c)) when "01101001101", 
		    std_logic_vector(to_unsigned(950, n_bits_c)) when "01101001110", 
		    std_logic_vector(to_unsigned(948, n_bits_c)) when "01101001111", 
		    std_logic_vector(to_unsigned(947, n_bits_c)) when "01101010000", 
		    std_logic_vector(to_unsigned(945, n_bits_c)) when "01101010001", 
		    std_logic_vector(to_unsigned(944, n_bits_c)) when "01101010010", 
		    std_logic_vector(to_unsigned(942, n_bits_c)) when "01101010011", 
		    std_logic_vector(to_unsigned(941, n_bits_c)) when "01101010100", 
		    std_logic_vector(to_unsigned(940, n_bits_c)) when "01101010101", 
		    std_logic_vector(to_unsigned(938, n_bits_c)) when "01101010110", 
		    std_logic_vector(to_unsigned(937, n_bits_c)) when "01101010111", 
		    std_logic_vector(to_unsigned(935, n_bits_c)) when "01101011000", 
		    std_logic_vector(to_unsigned(934, n_bits_c)) when "01101011001", 
		    std_logic_vector(to_unsigned(932, n_bits_c)) when "01101011010", 
		    std_logic_vector(to_unsigned(931, n_bits_c)) when "01101011011", 
		    std_logic_vector(to_unsigned(929, n_bits_c)) when "01101011100", 
		    std_logic_vector(to_unsigned(928, n_bits_c)) when "01101011101", 
		    std_logic_vector(to_unsigned(926, n_bits_c)) when "01101011110", 
		    std_logic_vector(to_unsigned(925, n_bits_c)) when "01101011111", 
		    std_logic_vector(to_unsigned(924, n_bits_c)) when "01101100000", 
		    std_logic_vector(to_unsigned(922, n_bits_c)) when "01101100001", 
		    std_logic_vector(to_unsigned(921, n_bits_c)) when "01101100010", 
		    std_logic_vector(to_unsigned(919, n_bits_c)) when "01101100011", 
		    std_logic_vector(to_unsigned(918, n_bits_c)) when "01101100100", 
		    std_logic_vector(to_unsigned(916, n_bits_c)) when "01101100101", 
		    std_logic_vector(to_unsigned(915, n_bits_c)) when "01101100110", 
		    std_logic_vector(to_unsigned(913, n_bits_c)) when "01101100111", 
		    std_logic_vector(to_unsigned(912, n_bits_c)) when "01101101000", 
		    std_logic_vector(to_unsigned(910, n_bits_c)) when "01101101001", 
		    std_logic_vector(to_unsigned(909, n_bits_c)) when "01101101010", 
		    std_logic_vector(to_unsigned(907, n_bits_c)) when "01101101011", 
		    std_logic_vector(to_unsigned(906, n_bits_c)) when "01101101100", 
		    std_logic_vector(to_unsigned(904, n_bits_c)) when "01101101101", 
		    std_logic_vector(to_unsigned(903, n_bits_c)) when "01101101110", 
		    std_logic_vector(to_unsigned(901, n_bits_c)) when "01101101111", 
		    std_logic_vector(to_unsigned(900, n_bits_c)) when "01101110000", 
		    std_logic_vector(to_unsigned(898, n_bits_c)) when "01101110001", 
		    std_logic_vector(to_unsigned(897, n_bits_c)) when "01101110010", 
		    std_logic_vector(to_unsigned(895, n_bits_c)) when "01101110011", 
		    std_logic_vector(to_unsigned(894, n_bits_c)) when "01101110100", 
		    std_logic_vector(to_unsigned(892, n_bits_c)) when "01101110101", 
		    std_logic_vector(to_unsigned(891, n_bits_c)) when "01101110110", 
		    std_logic_vector(to_unsigned(889, n_bits_c)) when "01101110111", 
		    std_logic_vector(to_unsigned(888, n_bits_c)) when "01101111000", 
		    std_logic_vector(to_unsigned(886, n_bits_c)) when "01101111001", 
		    std_logic_vector(to_unsigned(885, n_bits_c)) when "01101111010", 
		    std_logic_vector(to_unsigned(883, n_bits_c)) when "01101111011", 
		    std_logic_vector(to_unsigned(881, n_bits_c)) when "01101111100", 
		    std_logic_vector(to_unsigned(880, n_bits_c)) when "01101111101", 
		    std_logic_vector(to_unsigned(878, n_bits_c)) when "01101111110", 
		    std_logic_vector(to_unsigned(877, n_bits_c)) when "01101111111", 
		    std_logic_vector(to_unsigned(875, n_bits_c)) when "01110000000", 
		    std_logic_vector(to_unsigned(874, n_bits_c)) when "01110000001", 
		    std_logic_vector(to_unsigned(872, n_bits_c)) when "01110000010", 
		    std_logic_vector(to_unsigned(871, n_bits_c)) when "01110000011", 
		    std_logic_vector(to_unsigned(869, n_bits_c)) when "01110000100", 
		    std_logic_vector(to_unsigned(868, n_bits_c)) when "01110000101", 
		    std_logic_vector(to_unsigned(866, n_bits_c)) when "01110000110", 
		    std_logic_vector(to_unsigned(865, n_bits_c)) when "01110000111", 
		    std_logic_vector(to_unsigned(863, n_bits_c)) when "01110001000", 
		    std_logic_vector(to_unsigned(861, n_bits_c)) when "01110001001", 
		    std_logic_vector(to_unsigned(860, n_bits_c)) when "01110001010", 
		    std_logic_vector(to_unsigned(858, n_bits_c)) when "01110001011", 
		    std_logic_vector(to_unsigned(857, n_bits_c)) when "01110001100", 
		    std_logic_vector(to_unsigned(855, n_bits_c)) when "01110001101", 
		    std_logic_vector(to_unsigned(854, n_bits_c)) when "01110001110", 
		    std_logic_vector(to_unsigned(852, n_bits_c)) when "01110001111", 
		    std_logic_vector(to_unsigned(850, n_bits_c)) when "01110010000", 
		    std_logic_vector(to_unsigned(849, n_bits_c)) when "01110010001", 
		    std_logic_vector(to_unsigned(847, n_bits_c)) when "01110010010", 
		    std_logic_vector(to_unsigned(846, n_bits_c)) when "01110010011", 
		    std_logic_vector(to_unsigned(844, n_bits_c)) when "01110010100", 
		    std_logic_vector(to_unsigned(843, n_bits_c)) when "01110010101", 
		    std_logic_vector(to_unsigned(841, n_bits_c)) when "01110010110", 
		    std_logic_vector(to_unsigned(839, n_bits_c)) when "01110010111", 
		    std_logic_vector(to_unsigned(838, n_bits_c)) when "01110011000", 
		    std_logic_vector(to_unsigned(836, n_bits_c)) when "01110011001", 
		    std_logic_vector(to_unsigned(835, n_bits_c)) when "01110011010", 
		    std_logic_vector(to_unsigned(833, n_bits_c)) when "01110011011", 
		    std_logic_vector(to_unsigned(832, n_bits_c)) when "01110011100", 
		    std_logic_vector(to_unsigned(830, n_bits_c)) when "01110011101", 
		    std_logic_vector(to_unsigned(828, n_bits_c)) when "01110011110", 
		    std_logic_vector(to_unsigned(827, n_bits_c)) when "01110011111", 
		    std_logic_vector(to_unsigned(825, n_bits_c)) when "01110100000", 
		    std_logic_vector(to_unsigned(824, n_bits_c)) when "01110100001", 
		    std_logic_vector(to_unsigned(822, n_bits_c)) when "01110100010", 
		    std_logic_vector(to_unsigned(820, n_bits_c)) when "01110100011", 
		    std_logic_vector(to_unsigned(819, n_bits_c)) when "01110100100", 
		    std_logic_vector(to_unsigned(817, n_bits_c)) when "01110100101", 
		    std_logic_vector(to_unsigned(816, n_bits_c)) when "01110100110", 
		    std_logic_vector(to_unsigned(814, n_bits_c)) when "01110100111", 
		    std_logic_vector(to_unsigned(812, n_bits_c)) when "01110101000", 
		    std_logic_vector(to_unsigned(811, n_bits_c)) when "01110101001", 
		    std_logic_vector(to_unsigned(809, n_bits_c)) when "01110101010", 
		    std_logic_vector(to_unsigned(808, n_bits_c)) when "01110101011", 
		    std_logic_vector(to_unsigned(806, n_bits_c)) when "01110101100", 
		    std_logic_vector(to_unsigned(804, n_bits_c)) when "01110101101", 
		    std_logic_vector(to_unsigned(803, n_bits_c)) when "01110101110", 
		    std_logic_vector(to_unsigned(801, n_bits_c)) when "01110101111", 
		    std_logic_vector(to_unsigned(799, n_bits_c)) when "01110110000", 
		    std_logic_vector(to_unsigned(798, n_bits_c)) when "01110110001", 
		    std_logic_vector(to_unsigned(796, n_bits_c)) when "01110110010", 
		    std_logic_vector(to_unsigned(795, n_bits_c)) when "01110110011", 
		    std_logic_vector(to_unsigned(793, n_bits_c)) when "01110110100", 
		    std_logic_vector(to_unsigned(791, n_bits_c)) when "01110110101", 
		    std_logic_vector(to_unsigned(790, n_bits_c)) when "01110110110", 
		    std_logic_vector(to_unsigned(788, n_bits_c)) when "01110110111", 
		    std_logic_vector(to_unsigned(787, n_bits_c)) when "01110111000", 
		    std_logic_vector(to_unsigned(785, n_bits_c)) when "01110111001", 
		    std_logic_vector(to_unsigned(783, n_bits_c)) when "01110111010", 
		    std_logic_vector(to_unsigned(782, n_bits_c)) when "01110111011", 
		    std_logic_vector(to_unsigned(780, n_bits_c)) when "01110111100", 
		    std_logic_vector(to_unsigned(778, n_bits_c)) when "01110111101", 
		    std_logic_vector(to_unsigned(777, n_bits_c)) when "01110111110", 
		    std_logic_vector(to_unsigned(775, n_bits_c)) when "01110111111", 
		    std_logic_vector(to_unsigned(773, n_bits_c)) when "01111000000", 
		    std_logic_vector(to_unsigned(772, n_bits_c)) when "01111000001", 
		    std_logic_vector(to_unsigned(770, n_bits_c)) when "01111000010", 
		    std_logic_vector(to_unsigned(769, n_bits_c)) when "01111000011", 
		    std_logic_vector(to_unsigned(767, n_bits_c)) when "01111000100", 
		    std_logic_vector(to_unsigned(765, n_bits_c)) when "01111000101", 
		    std_logic_vector(to_unsigned(764, n_bits_c)) when "01111000110", 
		    std_logic_vector(to_unsigned(762, n_bits_c)) when "01111000111", 
		    std_logic_vector(to_unsigned(760, n_bits_c)) when "01111001000", 
		    std_logic_vector(to_unsigned(759, n_bits_c)) when "01111001001", 
		    std_logic_vector(to_unsigned(757, n_bits_c)) when "01111001010", 
		    std_logic_vector(to_unsigned(755, n_bits_c)) when "01111001011", 
		    std_logic_vector(to_unsigned(754, n_bits_c)) when "01111001100", 
		    std_logic_vector(to_unsigned(752, n_bits_c)) when "01111001101", 
		    std_logic_vector(to_unsigned(750, n_bits_c)) when "01111001110", 
		    std_logic_vector(to_unsigned(749, n_bits_c)) when "01111001111", 
		    std_logic_vector(to_unsigned(747, n_bits_c)) when "01111010000", 
		    std_logic_vector(to_unsigned(746, n_bits_c)) when "01111010001", 
		    std_logic_vector(to_unsigned(744, n_bits_c)) when "01111010010", 
		    std_logic_vector(to_unsigned(742, n_bits_c)) when "01111010011", 
		    std_logic_vector(to_unsigned(741, n_bits_c)) when "01111010100", 
		    std_logic_vector(to_unsigned(739, n_bits_c)) when "01111010101", 
		    std_logic_vector(to_unsigned(737, n_bits_c)) when "01111010110", 
		    std_logic_vector(to_unsigned(736, n_bits_c)) when "01111010111", 
		    std_logic_vector(to_unsigned(734, n_bits_c)) when "01111011000", 
		    std_logic_vector(to_unsigned(732, n_bits_c)) when "01111011001", 
		    std_logic_vector(to_unsigned(731, n_bits_c)) when "01111011010", 
		    std_logic_vector(to_unsigned(729, n_bits_c)) when "01111011011", 
		    std_logic_vector(to_unsigned(727, n_bits_c)) when "01111011100", 
		    std_logic_vector(to_unsigned(726, n_bits_c)) when "01111011101", 
		    std_logic_vector(to_unsigned(724, n_bits_c)) when "01111011110", 
		    std_logic_vector(to_unsigned(722, n_bits_c)) when "01111011111", 
		    std_logic_vector(to_unsigned(721, n_bits_c)) when "01111100000", 
		    std_logic_vector(to_unsigned(719, n_bits_c)) when "01111100001", 
		    std_logic_vector(to_unsigned(717, n_bits_c)) when "01111100010", 
		    std_logic_vector(to_unsigned(716, n_bits_c)) when "01111100011", 
		    std_logic_vector(to_unsigned(714, n_bits_c)) when "01111100100", 
		    std_logic_vector(to_unsigned(712, n_bits_c)) when "01111100101", 
		    std_logic_vector(to_unsigned(711, n_bits_c)) when "01111100110", 
		    std_logic_vector(to_unsigned(709, n_bits_c)) when "01111100111", 
		    std_logic_vector(to_unsigned(707, n_bits_c)) when "01111101000", 
		    std_logic_vector(to_unsigned(706, n_bits_c)) when "01111101001", 
		    std_logic_vector(to_unsigned(704, n_bits_c)) when "01111101010", 
		    std_logic_vector(to_unsigned(702, n_bits_c)) when "01111101011", 
		    std_logic_vector(to_unsigned(701, n_bits_c)) when "01111101100", 
		    std_logic_vector(to_unsigned(699, n_bits_c)) when "01111101101", 
		    std_logic_vector(to_unsigned(697, n_bits_c)) when "01111101110", 
		    std_logic_vector(to_unsigned(696, n_bits_c)) when "01111101111", 
		    std_logic_vector(to_unsigned(694, n_bits_c)) when "01111110000", 
		    std_logic_vector(to_unsigned(692, n_bits_c)) when "01111110001", 
		    std_logic_vector(to_unsigned(691, n_bits_c)) when "01111110010", 
		    std_logic_vector(to_unsigned(689, n_bits_c)) when "01111110011", 
		    std_logic_vector(to_unsigned(687, n_bits_c)) when "01111110100", 
		    std_logic_vector(to_unsigned(686, n_bits_c)) when "01111110101", 
		    std_logic_vector(to_unsigned(684, n_bits_c)) when "01111110110", 
		    std_logic_vector(to_unsigned(682, n_bits_c)) when "01111110111", 
		    std_logic_vector(to_unsigned(681, n_bits_c)) when "01111111000", 
		    std_logic_vector(to_unsigned(679, n_bits_c)) when "01111111001", 
		    std_logic_vector(to_unsigned(677, n_bits_c)) when "01111111010", 
		    std_logic_vector(to_unsigned(676, n_bits_c)) when "01111111011", 
		    std_logic_vector(to_unsigned(674, n_bits_c)) when "01111111100", 
		    std_logic_vector(to_unsigned(672, n_bits_c)) when "01111111101", 
		    std_logic_vector(to_unsigned(671, n_bits_c)) when "01111111110", 
		    std_logic_vector(to_unsigned(669, n_bits_c)) when "01111111111", 
		    std_logic_vector(to_unsigned(668, n_bits_c)) when "10000000000", 
		    std_logic_vector(to_unsigned(666, n_bits_c)) when "10000000001", 
		    std_logic_vector(to_unsigned(664, n_bits_c)) when "10000000010", 
		    std_logic_vector(to_unsigned(663, n_bits_c)) when "10000000011", 
		    std_logic_vector(to_unsigned(661, n_bits_c)) when "10000000100", 
		    std_logic_vector(to_unsigned(659, n_bits_c)) when "10000000101", 
		    std_logic_vector(to_unsigned(658, n_bits_c)) when "10000000110", 
		    std_logic_vector(to_unsigned(656, n_bits_c)) when "10000000111", 
		    std_logic_vector(to_unsigned(654, n_bits_c)) when "10000001000", 
		    std_logic_vector(to_unsigned(653, n_bits_c)) when "10000001001", 
		    std_logic_vector(to_unsigned(651, n_bits_c)) when "10000001010", 
		    std_logic_vector(to_unsigned(649, n_bits_c)) when "10000001011", 
		    std_logic_vector(to_unsigned(648, n_bits_c)) when "10000001100", 
		    std_logic_vector(to_unsigned(646, n_bits_c)) when "10000001101", 
		    std_logic_vector(to_unsigned(644, n_bits_c)) when "10000001110", 
		    std_logic_vector(to_unsigned(643, n_bits_c)) when "10000001111", 
		    std_logic_vector(to_unsigned(641, n_bits_c)) when "10000010000", 
		    std_logic_vector(to_unsigned(639, n_bits_c)) when "10000010001", 
		    std_logic_vector(to_unsigned(638, n_bits_c)) when "10000010010", 
		    std_logic_vector(to_unsigned(636, n_bits_c)) when "10000010011", 
		    std_logic_vector(to_unsigned(634, n_bits_c)) when "10000010100", 
		    std_logic_vector(to_unsigned(633, n_bits_c)) when "10000010101", 
		    std_logic_vector(to_unsigned(631, n_bits_c)) when "10000010110", 
		    std_logic_vector(to_unsigned(629, n_bits_c)) when "10000010111", 
		    std_logic_vector(to_unsigned(628, n_bits_c)) when "10000011000", 
		    std_logic_vector(to_unsigned(626, n_bits_c)) when "10000011001", 
		    std_logic_vector(to_unsigned(624, n_bits_c)) when "10000011010", 
		    std_logic_vector(to_unsigned(623, n_bits_c)) when "10000011011", 
		    std_logic_vector(to_unsigned(621, n_bits_c)) when "10000011100", 
		    std_logic_vector(to_unsigned(619, n_bits_c)) when "10000011101", 
		    std_logic_vector(to_unsigned(618, n_bits_c)) when "10000011110", 
		    std_logic_vector(to_unsigned(616, n_bits_c)) when "10000011111", 
		    std_logic_vector(to_unsigned(614, n_bits_c)) when "10000100000", 
		    std_logic_vector(to_unsigned(613, n_bits_c)) when "10000100001", 
		    std_logic_vector(to_unsigned(611, n_bits_c)) when "10000100010", 
		    std_logic_vector(to_unsigned(609, n_bits_c)) when "10000100011", 
		    std_logic_vector(to_unsigned(608, n_bits_c)) when "10000100100", 
		    std_logic_vector(to_unsigned(606, n_bits_c)) when "10000100101", 
		    std_logic_vector(to_unsigned(604, n_bits_c)) when "10000100110", 
		    std_logic_vector(to_unsigned(603, n_bits_c)) when "10000100111", 
		    std_logic_vector(to_unsigned(601, n_bits_c)) when "10000101000", 
		    std_logic_vector(to_unsigned(599, n_bits_c)) when "10000101001", 
		    std_logic_vector(to_unsigned(598, n_bits_c)) when "10000101010", 
		    std_logic_vector(to_unsigned(596, n_bits_c)) when "10000101011", 
		    std_logic_vector(to_unsigned(594, n_bits_c)) when "10000101100", 
		    std_logic_vector(to_unsigned(593, n_bits_c)) when "10000101101", 
		    std_logic_vector(to_unsigned(591, n_bits_c)) when "10000101110", 
		    std_logic_vector(to_unsigned(589, n_bits_c)) when "10000101111", 
		    std_logic_vector(to_unsigned(588, n_bits_c)) when "10000110000", 
		    std_logic_vector(to_unsigned(586, n_bits_c)) when "10000110001", 
		    std_logic_vector(to_unsigned(585, n_bits_c)) when "10000110010", 
		    std_logic_vector(to_unsigned(583, n_bits_c)) when "10000110011", 
		    std_logic_vector(to_unsigned(581, n_bits_c)) when "10000110100", 
		    std_logic_vector(to_unsigned(580, n_bits_c)) when "10000110101", 
		    std_logic_vector(to_unsigned(578, n_bits_c)) when "10000110110", 
		    std_logic_vector(to_unsigned(576, n_bits_c)) when "10000110111", 
		    std_logic_vector(to_unsigned(575, n_bits_c)) when "10000111000", 
		    std_logic_vector(to_unsigned(573, n_bits_c)) when "10000111001", 
		    std_logic_vector(to_unsigned(571, n_bits_c)) when "10000111010", 
		    std_logic_vector(to_unsigned(570, n_bits_c)) when "10000111011", 
		    std_logic_vector(to_unsigned(568, n_bits_c)) when "10000111100", 
		    std_logic_vector(to_unsigned(566, n_bits_c)) when "10000111101", 
		    std_logic_vector(to_unsigned(565, n_bits_c)) when "10000111110", 
		    std_logic_vector(to_unsigned(563, n_bits_c)) when "10000111111", 
		    std_logic_vector(to_unsigned(562, n_bits_c)) when "10001000000", 
		    std_logic_vector(to_unsigned(560, n_bits_c)) when "10001000001", 
		    std_logic_vector(to_unsigned(558, n_bits_c)) when "10001000010", 
		    std_logic_vector(to_unsigned(557, n_bits_c)) when "10001000011", 
		    std_logic_vector(to_unsigned(555, n_bits_c)) when "10001000100", 
		    std_logic_vector(to_unsigned(553, n_bits_c)) when "10001000101", 
		    std_logic_vector(to_unsigned(552, n_bits_c)) when "10001000110", 
		    std_logic_vector(to_unsigned(550, n_bits_c)) when "10001000111", 
		    std_logic_vector(to_unsigned(548, n_bits_c)) when "10001001000", 
		    std_logic_vector(to_unsigned(547, n_bits_c)) when "10001001001", 
		    std_logic_vector(to_unsigned(545, n_bits_c)) when "10001001010", 
		    std_logic_vector(to_unsigned(544, n_bits_c)) when "10001001011", 
		    std_logic_vector(to_unsigned(542, n_bits_c)) when "10001001100", 
		    std_logic_vector(to_unsigned(540, n_bits_c)) when "10001001101", 
		    std_logic_vector(to_unsigned(539, n_bits_c)) when "10001001110", 
		    std_logic_vector(to_unsigned(537, n_bits_c)) when "10001001111", 
		    std_logic_vector(to_unsigned(536, n_bits_c)) when "10001010000", 
		    std_logic_vector(to_unsigned(534, n_bits_c)) when "10001010001", 
		    std_logic_vector(to_unsigned(532, n_bits_c)) when "10001010010", 
		    std_logic_vector(to_unsigned(531, n_bits_c)) when "10001010011", 
		    std_logic_vector(to_unsigned(529, n_bits_c)) when "10001010100", 
		    std_logic_vector(to_unsigned(527, n_bits_c)) when "10001010101", 
		    std_logic_vector(to_unsigned(526, n_bits_c)) when "10001010110", 
		    std_logic_vector(to_unsigned(524, n_bits_c)) when "10001010111", 
		    std_logic_vector(to_unsigned(523, n_bits_c)) when "10001011000", 
		    std_logic_vector(to_unsigned(521, n_bits_c)) when "10001011001", 
		    std_logic_vector(to_unsigned(519, n_bits_c)) when "10001011010", 
		    std_logic_vector(to_unsigned(518, n_bits_c)) when "10001011011", 
		    std_logic_vector(to_unsigned(516, n_bits_c)) when "10001011100", 
		    std_logic_vector(to_unsigned(515, n_bits_c)) when "10001011101", 
		    std_logic_vector(to_unsigned(513, n_bits_c)) when "10001011110", 
		    std_logic_vector(to_unsigned(511, n_bits_c)) when "10001011111", 
		    std_logic_vector(to_unsigned(510, n_bits_c)) when "10001100000", 
		    std_logic_vector(to_unsigned(508, n_bits_c)) when "10001100001", 
		    std_logic_vector(to_unsigned(507, n_bits_c)) when "10001100010", 
		    std_logic_vector(to_unsigned(505, n_bits_c)) when "10001100011", 
		    std_logic_vector(to_unsigned(503, n_bits_c)) when "10001100100", 
		    std_logic_vector(to_unsigned(502, n_bits_c)) when "10001100101", 
		    std_logic_vector(to_unsigned(500, n_bits_c)) when "10001100110", 
		    std_logic_vector(to_unsigned(499, n_bits_c)) when "10001100111", 
		    std_logic_vector(to_unsigned(497, n_bits_c)) when "10001101000", 
		    std_logic_vector(to_unsigned(496, n_bits_c)) when "10001101001", 
		    std_logic_vector(to_unsigned(494, n_bits_c)) when "10001101010", 
		    std_logic_vector(to_unsigned(492, n_bits_c)) when "10001101011", 
		    std_logic_vector(to_unsigned(491, n_bits_c)) when "10001101100", 
		    std_logic_vector(to_unsigned(489, n_bits_c)) when "10001101101", 
		    std_logic_vector(to_unsigned(488, n_bits_c)) when "10001101110", 
		    std_logic_vector(to_unsigned(486, n_bits_c)) when "10001101111", 
		    std_logic_vector(to_unsigned(485, n_bits_c)) when "10001110000", 
		    std_logic_vector(to_unsigned(483, n_bits_c)) when "10001110001", 
		    std_logic_vector(to_unsigned(481, n_bits_c)) when "10001110010", 
		    std_logic_vector(to_unsigned(480, n_bits_c)) when "10001110011", 
		    std_logic_vector(to_unsigned(478, n_bits_c)) when "10001110100", 
		    std_logic_vector(to_unsigned(477, n_bits_c)) when "10001110101", 
		    std_logic_vector(to_unsigned(475, n_bits_c)) when "10001110110", 
		    std_logic_vector(to_unsigned(474, n_bits_c)) when "10001110111", 
		    std_logic_vector(to_unsigned(472, n_bits_c)) when "10001111000", 
		    std_logic_vector(to_unsigned(470, n_bits_c)) when "10001111001", 
		    std_logic_vector(to_unsigned(469, n_bits_c)) when "10001111010", 
		    std_logic_vector(to_unsigned(467, n_bits_c)) when "10001111011", 
		    std_logic_vector(to_unsigned(466, n_bits_c)) when "10001111100", 
		    std_logic_vector(to_unsigned(464, n_bits_c)) when "10001111101", 
		    std_logic_vector(to_unsigned(463, n_bits_c)) when "10001111110", 
		    std_logic_vector(to_unsigned(461, n_bits_c)) when "10001111111", 
		    std_logic_vector(to_unsigned(460, n_bits_c)) when "10010000000", 
		    std_logic_vector(to_unsigned(458, n_bits_c)) when "10010000001", 
		    std_logic_vector(to_unsigned(457, n_bits_c)) when "10010000010", 
		    std_logic_vector(to_unsigned(455, n_bits_c)) when "10010000011", 
		    std_logic_vector(to_unsigned(454, n_bits_c)) when "10010000100", 
		    std_logic_vector(to_unsigned(452, n_bits_c)) when "10010000101", 
		    std_logic_vector(to_unsigned(450, n_bits_c)) when "10010000110", 
		    std_logic_vector(to_unsigned(449, n_bits_c)) when "10010000111", 
		    std_logic_vector(to_unsigned(447, n_bits_c)) when "10010001000", 
		    std_logic_vector(to_unsigned(446, n_bits_c)) when "10010001001", 
		    std_logic_vector(to_unsigned(444, n_bits_c)) when "10010001010", 
		    std_logic_vector(to_unsigned(443, n_bits_c)) when "10010001011", 
		    std_logic_vector(to_unsigned(441, n_bits_c)) when "10010001100", 
		    std_logic_vector(to_unsigned(440, n_bits_c)) when "10010001101", 
		    std_logic_vector(to_unsigned(438, n_bits_c)) when "10010001110", 
		    std_logic_vector(to_unsigned(437, n_bits_c)) when "10010001111", 
		    std_logic_vector(to_unsigned(435, n_bits_c)) when "10010010000", 
		    std_logic_vector(to_unsigned(434, n_bits_c)) when "10010010001", 
		    std_logic_vector(to_unsigned(432, n_bits_c)) when "10010010010", 
		    std_logic_vector(to_unsigned(431, n_bits_c)) when "10010010011", 
		    std_logic_vector(to_unsigned(429, n_bits_c)) when "10010010100", 
		    std_logic_vector(to_unsigned(428, n_bits_c)) when "10010010101", 
		    std_logic_vector(to_unsigned(426, n_bits_c)) when "10010010110", 
		    std_logic_vector(to_unsigned(425, n_bits_c)) when "10010010111", 
		    std_logic_vector(to_unsigned(423, n_bits_c)) when "10010011000", 
		    std_logic_vector(to_unsigned(422, n_bits_c)) when "10010011001", 
		    std_logic_vector(to_unsigned(420, n_bits_c)) when "10010011010", 
		    std_logic_vector(to_unsigned(419, n_bits_c)) when "10010011011", 
		    std_logic_vector(to_unsigned(417, n_bits_c)) when "10010011100", 
		    std_logic_vector(to_unsigned(416, n_bits_c)) when "10010011101", 
		    std_logic_vector(to_unsigned(414, n_bits_c)) when "10010011110", 
		    std_logic_vector(to_unsigned(413, n_bits_c)) when "10010011111", 
		    std_logic_vector(to_unsigned(411, n_bits_c)) when "10010100000", 
		    std_logic_vector(to_unsigned(410, n_bits_c)) when "10010100001", 
		    std_logic_vector(to_unsigned(409, n_bits_c)) when "10010100010", 
		    std_logic_vector(to_unsigned(407, n_bits_c)) when "10010100011", 
		    std_logic_vector(to_unsigned(406, n_bits_c)) when "10010100100", 
		    std_logic_vector(to_unsigned(404, n_bits_c)) when "10010100101", 
		    std_logic_vector(to_unsigned(403, n_bits_c)) when "10010100110", 
		    std_logic_vector(to_unsigned(401, n_bits_c)) when "10010100111", 
		    std_logic_vector(to_unsigned(400, n_bits_c)) when "10010101000", 
		    std_logic_vector(to_unsigned(398, n_bits_c)) when "10010101001", 
		    std_logic_vector(to_unsigned(397, n_bits_c)) when "10010101010", 
		    std_logic_vector(to_unsigned(395, n_bits_c)) when "10010101011", 
		    std_logic_vector(to_unsigned(394, n_bits_c)) when "10010101100", 
		    std_logic_vector(to_unsigned(393, n_bits_c)) when "10010101101", 
		    std_logic_vector(to_unsigned(391, n_bits_c)) when "10010101110", 
		    std_logic_vector(to_unsigned(390, n_bits_c)) when "10010101111", 
		    std_logic_vector(to_unsigned(388, n_bits_c)) when "10010110000", 
		    std_logic_vector(to_unsigned(387, n_bits_c)) when "10010110001", 
		    std_logic_vector(to_unsigned(385, n_bits_c)) when "10010110010", 
		    std_logic_vector(to_unsigned(384, n_bits_c)) when "10010110011", 
		    std_logic_vector(to_unsigned(383, n_bits_c)) when "10010110100", 
		    std_logic_vector(to_unsigned(381, n_bits_c)) when "10010110101", 
		    std_logic_vector(to_unsigned(380, n_bits_c)) when "10010110110", 
		    std_logic_vector(to_unsigned(378, n_bits_c)) when "10010110111", 
		    std_logic_vector(to_unsigned(377, n_bits_c)) when "10010111000", 
		    std_logic_vector(to_unsigned(376, n_bits_c)) when "10010111001", 
		    std_logic_vector(to_unsigned(374, n_bits_c)) when "10010111010", 
		    std_logic_vector(to_unsigned(373, n_bits_c)) when "10010111011", 
		    std_logic_vector(to_unsigned(371, n_bits_c)) when "10010111100", 
		    std_logic_vector(to_unsigned(370, n_bits_c)) when "10010111101", 
		    std_logic_vector(to_unsigned(369, n_bits_c)) when "10010111110", 
		    std_logic_vector(to_unsigned(367, n_bits_c)) when "10010111111", 
		    std_logic_vector(to_unsigned(366, n_bits_c)) when "10011000000", 
		    std_logic_vector(to_unsigned(364, n_bits_c)) when "10011000001", 
		    std_logic_vector(to_unsigned(363, n_bits_c)) when "10011000010", 
		    std_logic_vector(to_unsigned(362, n_bits_c)) when "10011000011", 
		    std_logic_vector(to_unsigned(360, n_bits_c)) when "10011000100", 
		    std_logic_vector(to_unsigned(359, n_bits_c)) when "10011000101", 
		    std_logic_vector(to_unsigned(357, n_bits_c)) when "10011000110", 
		    std_logic_vector(to_unsigned(356, n_bits_c)) when "10011000111", 
		    std_logic_vector(to_unsigned(355, n_bits_c)) when "10011001000", 
		    std_logic_vector(to_unsigned(353, n_bits_c)) when "10011001001", 
		    std_logic_vector(to_unsigned(352, n_bits_c)) when "10011001010", 
		    std_logic_vector(to_unsigned(351, n_bits_c)) when "10011001011", 
		    std_logic_vector(to_unsigned(349, n_bits_c)) when "10011001100", 
		    std_logic_vector(to_unsigned(348, n_bits_c)) when "10011001101", 
		    std_logic_vector(to_unsigned(347, n_bits_c)) when "10011001110", 
		    std_logic_vector(to_unsigned(345, n_bits_c)) when "10011001111", 
		    std_logic_vector(to_unsigned(344, n_bits_c)) when "10011010000", 
		    std_logic_vector(to_unsigned(343, n_bits_c)) when "10011010001", 
		    std_logic_vector(to_unsigned(341, n_bits_c)) when "10011010010", 
		    std_logic_vector(to_unsigned(340, n_bits_c)) when "10011010011", 
		    std_logic_vector(to_unsigned(339, n_bits_c)) when "10011010100", 
		    std_logic_vector(to_unsigned(337, n_bits_c)) when "10011010101", 
		    std_logic_vector(to_unsigned(336, n_bits_c)) when "10011010110", 
		    std_logic_vector(to_unsigned(335, n_bits_c)) when "10011010111", 
		    std_logic_vector(to_unsigned(333, n_bits_c)) when "10011011000", 
		    std_logic_vector(to_unsigned(332, n_bits_c)) when "10011011001", 
		    std_logic_vector(to_unsigned(331, n_bits_c)) when "10011011010", 
		    std_logic_vector(to_unsigned(329, n_bits_c)) when "10011011011", 
		    std_logic_vector(to_unsigned(328, n_bits_c)) when "10011011100", 
		    std_logic_vector(to_unsigned(327, n_bits_c)) when "10011011101", 
		    std_logic_vector(to_unsigned(326, n_bits_c)) when "10011011110", 
		    std_logic_vector(to_unsigned(324, n_bits_c)) when "10011011111", 
		    std_logic_vector(to_unsigned(323, n_bits_c)) when "10011100000", 
		    std_logic_vector(to_unsigned(322, n_bits_c)) when "10011100001", 
		    std_logic_vector(to_unsigned(320, n_bits_c)) when "10011100010", 
		    std_logic_vector(to_unsigned(319, n_bits_c)) when "10011100011", 
		    std_logic_vector(to_unsigned(318, n_bits_c)) when "10011100100", 
		    std_logic_vector(to_unsigned(317, n_bits_c)) when "10011100101", 
		    std_logic_vector(to_unsigned(315, n_bits_c)) when "10011100110", 
		    std_logic_vector(to_unsigned(314, n_bits_c)) when "10011100111", 
		    std_logic_vector(to_unsigned(313, n_bits_c)) when "10011101000", 
		    std_logic_vector(to_unsigned(311, n_bits_c)) when "10011101001", 
		    std_logic_vector(to_unsigned(310, n_bits_c)) when "10011101010", 
		    std_logic_vector(to_unsigned(309, n_bits_c)) when "10011101011", 
		    std_logic_vector(to_unsigned(308, n_bits_c)) when "10011101100", 
		    std_logic_vector(to_unsigned(306, n_bits_c)) when "10011101101", 
		    std_logic_vector(to_unsigned(305, n_bits_c)) when "10011101110", 
		    std_logic_vector(to_unsigned(304, n_bits_c)) when "10011101111", 
		    std_logic_vector(to_unsigned(303, n_bits_c)) when "10011110000", 
		    std_logic_vector(to_unsigned(302, n_bits_c)) when "10011110001", 
		    std_logic_vector(to_unsigned(300, n_bits_c)) when "10011110010", 
		    std_logic_vector(to_unsigned(299, n_bits_c)) when "10011110011", 
		    std_logic_vector(to_unsigned(298, n_bits_c)) when "10011110100", 
		    std_logic_vector(to_unsigned(297, n_bits_c)) when "10011110101", 
		    std_logic_vector(to_unsigned(295, n_bits_c)) when "10011110110", 
		    std_logic_vector(to_unsigned(294, n_bits_c)) when "10011110111", 
		    std_logic_vector(to_unsigned(293, n_bits_c)) when "10011111000", 
		    std_logic_vector(to_unsigned(292, n_bits_c)) when "10011111001", 
		    std_logic_vector(to_unsigned(291, n_bits_c)) when "10011111010", 
		    std_logic_vector(to_unsigned(289, n_bits_c)) when "10011111011", 
		    std_logic_vector(to_unsigned(288, n_bits_c)) when "10011111100", 
		    std_logic_vector(to_unsigned(287, n_bits_c)) when "10011111101", 
		    std_logic_vector(to_unsigned(286, n_bits_c)) when "10011111110", 
		    std_logic_vector(to_unsigned(285, n_bits_c)) when "10011111111", 
		    std_logic_vector(to_unsigned(283, n_bits_c)) when "10100000000", 
		    std_logic_vector(to_unsigned(282, n_bits_c)) when "10100000001", 
		    std_logic_vector(to_unsigned(281, n_bits_c)) when "10100000010", 
		    std_logic_vector(to_unsigned(280, n_bits_c)) when "10100000011", 
		    std_logic_vector(to_unsigned(279, n_bits_c)) when "10100000100", 
		    std_logic_vector(to_unsigned(278, n_bits_c)) when "10100000101", 
		    std_logic_vector(to_unsigned(276, n_bits_c)) when "10100000110", 
		    std_logic_vector(to_unsigned(275, n_bits_c)) when "10100000111", 
		    std_logic_vector(to_unsigned(274, n_bits_c)) when "10100001000", 
		    std_logic_vector(to_unsigned(273, n_bits_c)) when "10100001001", 
		    std_logic_vector(to_unsigned(272, n_bits_c)) when "10100001010", 
		    std_logic_vector(to_unsigned(271, n_bits_c)) when "10100001011", 
		    std_logic_vector(to_unsigned(270, n_bits_c)) when "10100001100", 
		    std_logic_vector(to_unsigned(268, n_bits_c)) when "10100001101", 
		    std_logic_vector(to_unsigned(267, n_bits_c)) when "10100001110", 
		    std_logic_vector(to_unsigned(266, n_bits_c)) when "10100001111", 
		    std_logic_vector(to_unsigned(265, n_bits_c)) when "10100010000", 
		    std_logic_vector(to_unsigned(264, n_bits_c)) when "10100010001", 
		    std_logic_vector(to_unsigned(263, n_bits_c)) when "10100010010", 
		    std_logic_vector(to_unsigned(262, n_bits_c)) when "10100010011", 
		    std_logic_vector(to_unsigned(261, n_bits_c)) when "10100010100", 
		    std_logic_vector(to_unsigned(260, n_bits_c)) when "10100010101", 
		    std_logic_vector(to_unsigned(258, n_bits_c)) when "10100010110", 
		    std_logic_vector(to_unsigned(257, n_bits_c)) when "10100010111", 
		    std_logic_vector(to_unsigned(256, n_bits_c)) when "10100011000", 
		    std_logic_vector(to_unsigned(255, n_bits_c)) when "10100011001", 
		    std_logic_vector(to_unsigned(254, n_bits_c)) when "10100011010", 
		    std_logic_vector(to_unsigned(253, n_bits_c)) when "10100011011", 
		    std_logic_vector(to_unsigned(252, n_bits_c)) when "10100011100", 
		    std_logic_vector(to_unsigned(251, n_bits_c)) when "10100011101", 
		    std_logic_vector(to_unsigned(250, n_bits_c)) when "10100011110", 
		    std_logic_vector(to_unsigned(249, n_bits_c)) when "10100011111", 
		    std_logic_vector(to_unsigned(248, n_bits_c)) when "10100100000", 
		    std_logic_vector(to_unsigned(247, n_bits_c)) when "10100100001", 
		    std_logic_vector(to_unsigned(246, n_bits_c)) when "10100100010", 
		    std_logic_vector(to_unsigned(244, n_bits_c)) when "10100100011", 
		    std_logic_vector(to_unsigned(243, n_bits_c)) when "10100100100", 
		    std_logic_vector(to_unsigned(242, n_bits_c)) when "10100100101", 
		    std_logic_vector(to_unsigned(241, n_bits_c)) when "10100100110", 
		    std_logic_vector(to_unsigned(240, n_bits_c)) when "10100100111", 
		    std_logic_vector(to_unsigned(239, n_bits_c)) when "10100101000", 
		    std_logic_vector(to_unsigned(238, n_bits_c)) when "10100101001", 
		    std_logic_vector(to_unsigned(237, n_bits_c)) when "10100101010", 
		    std_logic_vector(to_unsigned(236, n_bits_c)) when "10100101011", 
		    std_logic_vector(to_unsigned(235, n_bits_c)) when "10100101100", 
		    std_logic_vector(to_unsigned(234, n_bits_c)) when "10100101101", 
		    std_logic_vector(to_unsigned(233, n_bits_c)) when "10100101110", 
		    std_logic_vector(to_unsigned(232, n_bits_c)) when "10100101111", 
		    std_logic_vector(to_unsigned(231, n_bits_c)) when "10100110000", 
		    std_logic_vector(to_unsigned(230, n_bits_c)) when "10100110001", 
		    std_logic_vector(to_unsigned(229, n_bits_c)) when "10100110010", 
		    std_logic_vector(to_unsigned(228, n_bits_c)) when "10100110011", 
		    std_logic_vector(to_unsigned(227, n_bits_c)) when "10100110100", 
		    std_logic_vector(to_unsigned(226, n_bits_c)) when "10100110101", 
		    std_logic_vector(to_unsigned(225, n_bits_c)) when "10100110110", 
		    std_logic_vector(to_unsigned(224, n_bits_c)) when "10100110111", 
		    std_logic_vector(to_unsigned(223, n_bits_c)) when "10100111000", 
		    std_logic_vector(to_unsigned(222, n_bits_c)) when "10100111001", 
		    std_logic_vector(to_unsigned(222, n_bits_c)) when "10100111010", 
		    std_logic_vector(to_unsigned(221, n_bits_c)) when "10100111011", 
		    std_logic_vector(to_unsigned(220, n_bits_c)) when "10100111100", 
		    std_logic_vector(to_unsigned(219, n_bits_c)) when "10100111101", 
		    std_logic_vector(to_unsigned(218, n_bits_c)) when "10100111110", 
		    std_logic_vector(to_unsigned(217, n_bits_c)) when "10100111111", 
		    std_logic_vector(to_unsigned(216, n_bits_c)) when "10101000000", 
		    std_logic_vector(to_unsigned(215, n_bits_c)) when "10101000001", 
		    std_logic_vector(to_unsigned(214, n_bits_c)) when "10101000010", 
		    std_logic_vector(to_unsigned(213, n_bits_c)) when "10101000011", 
		    std_logic_vector(to_unsigned(212, n_bits_c)) when "10101000100", 
		    std_logic_vector(to_unsigned(211, n_bits_c)) when "10101000101", 
		    std_logic_vector(to_unsigned(210, n_bits_c)) when "10101000110", 
		    std_logic_vector(to_unsigned(210, n_bits_c)) when "10101000111", 
		    std_logic_vector(to_unsigned(209, n_bits_c)) when "10101001000", 
		    std_logic_vector(to_unsigned(208, n_bits_c)) when "10101001001", 
		    std_logic_vector(to_unsigned(207, n_bits_c)) when "10101001010", 
		    std_logic_vector(to_unsigned(206, n_bits_c)) when "10101001011", 
		    std_logic_vector(to_unsigned(205, n_bits_c)) when "10101001100", 
		    std_logic_vector(to_unsigned(204, n_bits_c)) when "10101001101", 
		    std_logic_vector(to_unsigned(203, n_bits_c)) when "10101001110", 
		    std_logic_vector(to_unsigned(202, n_bits_c)) when "10101001111", 
		    std_logic_vector(to_unsigned(202, n_bits_c)) when "10101010000", 
		    std_logic_vector(to_unsigned(201, n_bits_c)) when "10101010001", 
		    std_logic_vector(to_unsigned(200, n_bits_c)) when "10101010010", 
		    std_logic_vector(to_unsigned(199, n_bits_c)) when "10101010011", 
		    std_logic_vector(to_unsigned(198, n_bits_c)) when "10101010100", 
		    std_logic_vector(to_unsigned(197, n_bits_c)) when "10101010101", 
		    std_logic_vector(to_unsigned(197, n_bits_c)) when "10101010110", 
		    std_logic_vector(to_unsigned(196, n_bits_c)) when "10101010111", 
		    std_logic_vector(to_unsigned(195, n_bits_c)) when "10101011000", 
		    std_logic_vector(to_unsigned(194, n_bits_c)) when "10101011001", 
		    std_logic_vector(to_unsigned(193, n_bits_c)) when "10101011010", 
		    std_logic_vector(to_unsigned(192, n_bits_c)) when "10101011011", 
		    std_logic_vector(to_unsigned(192, n_bits_c)) when "10101011100", 
		    std_logic_vector(to_unsigned(191, n_bits_c)) when "10101011101", 
		    std_logic_vector(to_unsigned(190, n_bits_c)) when "10101011110", 
		    std_logic_vector(to_unsigned(189, n_bits_c)) when "10101011111", 
		    std_logic_vector(to_unsigned(188, n_bits_c)) when "10101100000", 
		    std_logic_vector(to_unsigned(188, n_bits_c)) when "10101100001", 
		    std_logic_vector(to_unsigned(187, n_bits_c)) when "10101100010", 
		    std_logic_vector(to_unsigned(186, n_bits_c)) when "10101100011", 
		    std_logic_vector(to_unsigned(185, n_bits_c)) when "10101100100", 
		    std_logic_vector(to_unsigned(185, n_bits_c)) when "10101100101", 
		    std_logic_vector(to_unsigned(184, n_bits_c)) when "10101100110", 
		    std_logic_vector(to_unsigned(183, n_bits_c)) when "10101100111", 
		    std_logic_vector(to_unsigned(182, n_bits_c)) when "10101101000", 
		    std_logic_vector(to_unsigned(182, n_bits_c)) when "10101101001", 
		    std_logic_vector(to_unsigned(181, n_bits_c)) when "10101101010", 
		    std_logic_vector(to_unsigned(180, n_bits_c)) when "10101101011", 
		    std_logic_vector(to_unsigned(179, n_bits_c)) when "10101101100", 
		    std_logic_vector(to_unsigned(179, n_bits_c)) when "10101101101", 
		    std_logic_vector(to_unsigned(178, n_bits_c)) when "10101101110", 
		    std_logic_vector(to_unsigned(177, n_bits_c)) when "10101101111", 
		    std_logic_vector(to_unsigned(177, n_bits_c)) when "10101110000", 
		    std_logic_vector(to_unsigned(176, n_bits_c)) when "10101110001", 
		    std_logic_vector(to_unsigned(175, n_bits_c)) when "10101110010", 
		    std_logic_vector(to_unsigned(174, n_bits_c)) when "10101110011", 
		    std_logic_vector(to_unsigned(174, n_bits_c)) when "10101110100", 
		    std_logic_vector(to_unsigned(173, n_bits_c)) when "10101110101", 
		    std_logic_vector(to_unsigned(172, n_bits_c)) when "10101110110", 
		    std_logic_vector(to_unsigned(172, n_bits_c)) when "10101110111", 
		    std_logic_vector(to_unsigned(171, n_bits_c)) when "10101111000", 
		    std_logic_vector(to_unsigned(170, n_bits_c)) when "10101111001", 
		    std_logic_vector(to_unsigned(170, n_bits_c)) when "10101111010", 
		    std_logic_vector(to_unsigned(169, n_bits_c)) when "10101111011", 
		    std_logic_vector(to_unsigned(168, n_bits_c)) when "10101111100", 
		    std_logic_vector(to_unsigned(168, n_bits_c)) when "10101111101", 
		    std_logic_vector(to_unsigned(167, n_bits_c)) when "10101111110", 
		    std_logic_vector(to_unsigned(166, n_bits_c)) when "10101111111", 
		    std_logic_vector(to_unsigned(166, n_bits_c)) when "10110000000", 
		    std_logic_vector(to_unsigned(165, n_bits_c)) when "10110000001", 
		    std_logic_vector(to_unsigned(164, n_bits_c)) when "10110000010", 
		    std_logic_vector(to_unsigned(164, n_bits_c)) when "10110000011", 
		    std_logic_vector(to_unsigned(163, n_bits_c)) when "10110000100", 
		    std_logic_vector(to_unsigned(163, n_bits_c)) when "10110000101", 
		    std_logic_vector(to_unsigned(162, n_bits_c)) when "10110000110", 
		    std_logic_vector(to_unsigned(161, n_bits_c)) when "10110000111", 
		    std_logic_vector(to_unsigned(161, n_bits_c)) when "10110001000", 
		    std_logic_vector(to_unsigned(160, n_bits_c)) when "10110001001", 
		    std_logic_vector(to_unsigned(160, n_bits_c)) when "10110001010", 
		    std_logic_vector(to_unsigned(159, n_bits_c)) when "10110001011", 
		    std_logic_vector(to_unsigned(158, n_bits_c)) when "10110001100", 
		    std_logic_vector(to_unsigned(158, n_bits_c)) when "10110001101", 
		    std_logic_vector(to_unsigned(157, n_bits_c)) when "10110001110", 
		    std_logic_vector(to_unsigned(157, n_bits_c)) when "10110001111", 
		    std_logic_vector(to_unsigned(156, n_bits_c)) when "10110010000", 
		    std_logic_vector(to_unsigned(156, n_bits_c)) when "10110010001", 
		    std_logic_vector(to_unsigned(155, n_bits_c)) when "10110010010", 
		    std_logic_vector(to_unsigned(154, n_bits_c)) when "10110010011", 
		    std_logic_vector(to_unsigned(154, n_bits_c)) when "10110010100", 
		    std_logic_vector(to_unsigned(153, n_bits_c)) when "10110010101", 
		    std_logic_vector(to_unsigned(153, n_bits_c)) when "10110010110", 
		    std_logic_vector(to_unsigned(152, n_bits_c)) when "10110010111", 
		    std_logic_vector(to_unsigned(152, n_bits_c)) when "10110011000", 
		    std_logic_vector(to_unsigned(151, n_bits_c)) when "10110011001", 
		    std_logic_vector(to_unsigned(151, n_bits_c)) when "10110011010", 
		    std_logic_vector(to_unsigned(150, n_bits_c)) when "10110011011", 
		    std_logic_vector(to_unsigned(150, n_bits_c)) when "10110011100", 
		    std_logic_vector(to_unsigned(149, n_bits_c)) when "10110011101", 
		    std_logic_vector(to_unsigned(149, n_bits_c)) when "10110011110", 
		    std_logic_vector(to_unsigned(148, n_bits_c)) when "10110011111", 
		    std_logic_vector(to_unsigned(148, n_bits_c)) when "10110100000", 
		    std_logic_vector(to_unsigned(147, n_bits_c)) when "10110100001", 
		    std_logic_vector(to_unsigned(147, n_bits_c)) when "10110100010", 
		    std_logic_vector(to_unsigned(146, n_bits_c)) when "10110100011", 
		    std_logic_vector(to_unsigned(146, n_bits_c)) when "10110100100", 
		    std_logic_vector(to_unsigned(145, n_bits_c)) when "10110100101", 
		    std_logic_vector(to_unsigned(145, n_bits_c)) when "10110100110", 
		    std_logic_vector(to_unsigned(144, n_bits_c)) when "10110100111", 
		    std_logic_vector(to_unsigned(144, n_bits_c)) when "10110101000", 
		    std_logic_vector(to_unsigned(144, n_bits_c)) when "10110101001", 
		    std_logic_vector(to_unsigned(143, n_bits_c)) when "10110101010", 
		    std_logic_vector(to_unsigned(143, n_bits_c)) when "10110101011", 
		    std_logic_vector(to_unsigned(142, n_bits_c)) when "10110101100", 
		    std_logic_vector(to_unsigned(142, n_bits_c)) when "10110101101", 
		    std_logic_vector(to_unsigned(141, n_bits_c)) when "10110101110", 
		    std_logic_vector(to_unsigned(141, n_bits_c)) when "10110101111", 
		    std_logic_vector(to_unsigned(141, n_bits_c)) when "10110110000", 
		    std_logic_vector(to_unsigned(140, n_bits_c)) when "10110110001", 
		    std_logic_vector(to_unsigned(140, n_bits_c)) when "10110110010", 
		    std_logic_vector(to_unsigned(139, n_bits_c)) when "10110110011", 
		    std_logic_vector(to_unsigned(139, n_bits_c)) when "10110110100", 
		    std_logic_vector(to_unsigned(139, n_bits_c)) when "10110110101", 
		    std_logic_vector(to_unsigned(138, n_bits_c)) when "10110110110", 
		    std_logic_vector(to_unsigned(138, n_bits_c)) when "10110110111", 
		    std_logic_vector(to_unsigned(138, n_bits_c)) when "10110111000", 
		    std_logic_vector(to_unsigned(137, n_bits_c)) when "10110111001", 
		    std_logic_vector(to_unsigned(137, n_bits_c)) when "10110111010", 
		    std_logic_vector(to_unsigned(136, n_bits_c)) when "10110111011", 
		    std_logic_vector(to_unsigned(136, n_bits_c)) when "10110111100", 
		    std_logic_vector(to_unsigned(136, n_bits_c)) when "10110111101", 
		    std_logic_vector(to_unsigned(135, n_bits_c)) when "10110111110", 
		    std_logic_vector(to_unsigned(135, n_bits_c)) when "10110111111", 
		    std_logic_vector(to_unsigned(135, n_bits_c)) when "10111000000", 
		    std_logic_vector(to_unsigned(134, n_bits_c)) when "10111000001", 
		    std_logic_vector(to_unsigned(134, n_bits_c)) when "10111000010", 
		    std_logic_vector(to_unsigned(134, n_bits_c)) when "10111000011", 
		    std_logic_vector(to_unsigned(134, n_bits_c)) when "10111000100", 
		    std_logic_vector(to_unsigned(133, n_bits_c)) when "10111000101", 
		    std_logic_vector(to_unsigned(133, n_bits_c)) when "10111000110", 
		    std_logic_vector(to_unsigned(133, n_bits_c)) when "10111000111", 
		    std_logic_vector(to_unsigned(132, n_bits_c)) when "10111001000", 
		    std_logic_vector(to_unsigned(132, n_bits_c)) when "10111001001", 
		    std_logic_vector(to_unsigned(132, n_bits_c)) when "10111001010", 
		    std_logic_vector(to_unsigned(132, n_bits_c)) when "10111001011", 
		    std_logic_vector(to_unsigned(131, n_bits_c)) when "10111001100", 
		    std_logic_vector(to_unsigned(131, n_bits_c)) when "10111001101", 
		    std_logic_vector(to_unsigned(131, n_bits_c)) when "10111001110", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "10111001111", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "10111010000", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "10111010001", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "10111010010", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "10111010011", 
		    std_logic_vector(to_unsigned(129, n_bits_c)) when "10111010100", 
		    std_logic_vector(to_unsigned(129, n_bits_c)) when "10111010101", 
		    std_logic_vector(to_unsigned(129, n_bits_c)) when "10111010110", 
		    std_logic_vector(to_unsigned(129, n_bits_c)) when "10111010111", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "10111011000", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "10111011001", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "10111011010", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "10111011011", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "10111011100", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "10111011101", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "10111011110", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "10111011111", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "10111100000", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "10111100001", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "10111100010", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "10111100011", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "10111100100", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "10111100101", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "10111100110", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "10111100111", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "10111101000", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "10111101001", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "10111101010", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111101011", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111101100", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111101101", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111101110", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111101111", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111110000", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111110001", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111110010", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111110011", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111110100", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111110101", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111110110", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111110111", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "10111111000", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "10111111001", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "10111111010", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "10111111011", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "10111111100", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "10111111101", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "10111111110", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "10111111111", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "11000000000", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "11000000001", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "11000000010", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "11000000011", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "11000000100", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "11000000101", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "11000000110", 
		    std_logic_vector(to_unsigned(124, n_bits_c)) when "11000000111", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000001000", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000001001", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000001010", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000001011", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000001100", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000001101", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000001110", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000001111", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000010000", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000010001", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000010010", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000010011", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000010100", 
		    std_logic_vector(to_unsigned(125, n_bits_c)) when "11000010101", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "11000010110", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "11000010111", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "11000011000", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "11000011001", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "11000011010", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "11000011011", 
		    std_logic_vector(to_unsigned(126, n_bits_c)) when "11000011100", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "11000011101", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "11000011110", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "11000011111", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "11000100000", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "11000100001", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "11000100010", 
		    std_logic_vector(to_unsigned(127, n_bits_c)) when "11000100011", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "11000100100", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "11000100101", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "11000100110", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "11000100111", 
		    std_logic_vector(to_unsigned(128, n_bits_c)) when "11000101000", 
		    std_logic_vector(to_unsigned(129, n_bits_c)) when "11000101001", 
		    std_logic_vector(to_unsigned(129, n_bits_c)) when "11000101010", 
		    std_logic_vector(to_unsigned(129, n_bits_c)) when "11000101011", 
		    std_logic_vector(to_unsigned(129, n_bits_c)) when "11000101100", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "11000101101", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "11000101110", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "11000101111", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "11000110000", 
		    std_logic_vector(to_unsigned(130, n_bits_c)) when "11000110001", 
		    std_logic_vector(to_unsigned(131, n_bits_c)) when "11000110010", 
		    std_logic_vector(to_unsigned(131, n_bits_c)) when "11000110011", 
		    std_logic_vector(to_unsigned(131, n_bits_c)) when "11000110100", 
		    std_logic_vector(to_unsigned(132, n_bits_c)) when "11000110101", 
		    std_logic_vector(to_unsigned(132, n_bits_c)) when "11000110110", 
		    std_logic_vector(to_unsigned(132, n_bits_c)) when "11000110111", 
		    std_logic_vector(to_unsigned(132, n_bits_c)) when "11000111000", 
		    std_logic_vector(to_unsigned(133, n_bits_c)) when "11000111001", 
		    std_logic_vector(to_unsigned(133, n_bits_c)) when "11000111010", 
		    std_logic_vector(to_unsigned(133, n_bits_c)) when "11000111011", 
		    std_logic_vector(to_unsigned(134, n_bits_c)) when "11000111100", 
		    std_logic_vector(to_unsigned(134, n_bits_c)) when "11000111101", 
		    std_logic_vector(to_unsigned(134, n_bits_c)) when "11000111110", 
		    std_logic_vector(to_unsigned(134, n_bits_c)) when "11000111111", 
		    std_logic_vector(to_unsigned(135, n_bits_c)) when "11001000000", 
		    std_logic_vector(to_unsigned(135, n_bits_c)) when "11001000001", 
		    std_logic_vector(to_unsigned(135, n_bits_c)) when "11001000010", 
		    std_logic_vector(to_unsigned(136, n_bits_c)) when "11001000011", 
		    std_logic_vector(to_unsigned(136, n_bits_c)) when "11001000100", 
		    std_logic_vector(to_unsigned(136, n_bits_c)) when "11001000101", 
		    std_logic_vector(to_unsigned(137, n_bits_c)) when "11001000110", 
		    std_logic_vector(to_unsigned(137, n_bits_c)) when "11001000111", 
		    std_logic_vector(to_unsigned(138, n_bits_c)) when "11001001000", 
		    std_logic_vector(to_unsigned(138, n_bits_c)) when "11001001001", 
		    std_logic_vector(to_unsigned(138, n_bits_c)) when "11001001010", 
		    std_logic_vector(to_unsigned(139, n_bits_c)) when "11001001011", 
		    std_logic_vector(to_unsigned(139, n_bits_c)) when "11001001100", 
		    std_logic_vector(to_unsigned(139, n_bits_c)) when "11001001101", 
		    std_logic_vector(to_unsigned(140, n_bits_c)) when "11001001110", 
		    std_logic_vector(to_unsigned(140, n_bits_c)) when "11001001111", 
		    std_logic_vector(to_unsigned(141, n_bits_c)) when "11001010000", 
		    std_logic_vector(to_unsigned(141, n_bits_c)) when "11001010001", 
		    std_logic_vector(to_unsigned(141, n_bits_c)) when "11001010010", 
		    std_logic_vector(to_unsigned(142, n_bits_c)) when "11001010011", 
		    std_logic_vector(to_unsigned(142, n_bits_c)) when "11001010100", 
		    std_logic_vector(to_unsigned(143, n_bits_c)) when "11001010101", 
		    std_logic_vector(to_unsigned(143, n_bits_c)) when "11001010110", 
		    std_logic_vector(to_unsigned(144, n_bits_c)) when "11001010111", 
		    std_logic_vector(to_unsigned(144, n_bits_c)) when "11001011000", 
		    std_logic_vector(to_unsigned(144, n_bits_c)) when "11001011001", 
		    std_logic_vector(to_unsigned(145, n_bits_c)) when "11001011010", 
		    std_logic_vector(to_unsigned(145, n_bits_c)) when "11001011011", 
		    std_logic_vector(to_unsigned(146, n_bits_c)) when "11001011100", 
		    std_logic_vector(to_unsigned(146, n_bits_c)) when "11001011101", 
		    std_logic_vector(to_unsigned(147, n_bits_c)) when "11001011110", 
		    std_logic_vector(to_unsigned(147, n_bits_c)) when "11001011111", 
		    std_logic_vector(to_unsigned(148, n_bits_c)) when "11001100000", 
		    std_logic_vector(to_unsigned(148, n_bits_c)) when "11001100001", 
		    std_logic_vector(to_unsigned(149, n_bits_c)) when "11001100010", 
		    std_logic_vector(to_unsigned(149, n_bits_c)) when "11001100011", 
		    std_logic_vector(to_unsigned(150, n_bits_c)) when "11001100100", 
		    std_logic_vector(to_unsigned(150, n_bits_c)) when "11001100101", 
		    std_logic_vector(to_unsigned(151, n_bits_c)) when "11001100110", 
		    std_logic_vector(to_unsigned(151, n_bits_c)) when "11001100111", 
		    std_logic_vector(to_unsigned(152, n_bits_c)) when "11001101000", 
		    std_logic_vector(to_unsigned(152, n_bits_c)) when "11001101001", 
		    std_logic_vector(to_unsigned(153, n_bits_c)) when "11001101010", 
		    std_logic_vector(to_unsigned(153, n_bits_c)) when "11001101011", 
		    std_logic_vector(to_unsigned(154, n_bits_c)) when "11001101100", 
		    std_logic_vector(to_unsigned(154, n_bits_c)) when "11001101101", 
		    std_logic_vector(to_unsigned(155, n_bits_c)) when "11001101110", 
		    std_logic_vector(to_unsigned(156, n_bits_c)) when "11001101111", 
		    std_logic_vector(to_unsigned(156, n_bits_c)) when "11001110000", 
		    std_logic_vector(to_unsigned(157, n_bits_c)) when "11001110001", 
		    std_logic_vector(to_unsigned(157, n_bits_c)) when "11001110010", 
		    std_logic_vector(to_unsigned(158, n_bits_c)) when "11001110011", 
		    std_logic_vector(to_unsigned(158, n_bits_c)) when "11001110100", 
		    std_logic_vector(to_unsigned(159, n_bits_c)) when "11001110101", 
		    std_logic_vector(to_unsigned(160, n_bits_c)) when "11001110110", 
		    std_logic_vector(to_unsigned(160, n_bits_c)) when "11001110111", 
		    std_logic_vector(to_unsigned(161, n_bits_c)) when "11001111000", 
		    std_logic_vector(to_unsigned(161, n_bits_c)) when "11001111001", 
		    std_logic_vector(to_unsigned(162, n_bits_c)) when "11001111010", 
		    std_logic_vector(to_unsigned(163, n_bits_c)) when "11001111011", 
		    std_logic_vector(to_unsigned(163, n_bits_c)) when "11001111100", 
		    std_logic_vector(to_unsigned(164, n_bits_c)) when "11001111101", 
		    std_logic_vector(to_unsigned(164, n_bits_c)) when "11001111110", 
		    std_logic_vector(to_unsigned(165, n_bits_c)) when "11001111111", 
		    std_logic_vector(to_unsigned(166, n_bits_c)) when "11010000000", 
		    std_logic_vector(to_unsigned(166, n_bits_c)) when "11010000001", 
		    std_logic_vector(to_unsigned(167, n_bits_c)) when "11010000010", 
		    std_logic_vector(to_unsigned(168, n_bits_c)) when "11010000011", 
		    std_logic_vector(to_unsigned(168, n_bits_c)) when "11010000100", 
		    std_logic_vector(to_unsigned(169, n_bits_c)) when "11010000101", 
		    std_logic_vector(to_unsigned(170, n_bits_c)) when "11010000110", 
		    std_logic_vector(to_unsigned(170, n_bits_c)) when "11010000111", 
		    std_logic_vector(to_unsigned(171, n_bits_c)) when "11010001000", 
		    std_logic_vector(to_unsigned(172, n_bits_c)) when "11010001001", 
		    std_logic_vector(to_unsigned(172, n_bits_c)) when "11010001010", 
		    std_logic_vector(to_unsigned(173, n_bits_c)) when "11010001011", 
		    std_logic_vector(to_unsigned(174, n_bits_c)) when "11010001100", 
		    std_logic_vector(to_unsigned(174, n_bits_c)) when "11010001101", 
		    std_logic_vector(to_unsigned(175, n_bits_c)) when "11010001110", 
		    std_logic_vector(to_unsigned(176, n_bits_c)) when "11010001111", 
		    std_logic_vector(to_unsigned(177, n_bits_c)) when "11010010000", 
		    std_logic_vector(to_unsigned(177, n_bits_c)) when "11010010001", 
		    std_logic_vector(to_unsigned(178, n_bits_c)) when "11010010010", 
		    std_logic_vector(to_unsigned(179, n_bits_c)) when "11010010011", 
		    std_logic_vector(to_unsigned(179, n_bits_c)) when "11010010100", 
		    std_logic_vector(to_unsigned(180, n_bits_c)) when "11010010101", 
		    std_logic_vector(to_unsigned(181, n_bits_c)) when "11010010110", 
		    std_logic_vector(to_unsigned(182, n_bits_c)) when "11010010111", 
		    std_logic_vector(to_unsigned(182, n_bits_c)) when "11010011000", 
		    std_logic_vector(to_unsigned(183, n_bits_c)) when "11010011001", 
		    std_logic_vector(to_unsigned(184, n_bits_c)) when "11010011010", 
		    std_logic_vector(to_unsigned(185, n_bits_c)) when "11010011011", 
		    std_logic_vector(to_unsigned(185, n_bits_c)) when "11010011100", 
		    std_logic_vector(to_unsigned(186, n_bits_c)) when "11010011101", 
		    std_logic_vector(to_unsigned(187, n_bits_c)) when "11010011110", 
		    std_logic_vector(to_unsigned(188, n_bits_c)) when "11010011111", 
		    std_logic_vector(to_unsigned(188, n_bits_c)) when "11010100000", 
		    std_logic_vector(to_unsigned(189, n_bits_c)) when "11010100001", 
		    std_logic_vector(to_unsigned(190, n_bits_c)) when "11010100010", 
		    std_logic_vector(to_unsigned(191, n_bits_c)) when "11010100011", 
		    std_logic_vector(to_unsigned(192, n_bits_c)) when "11010100100", 
		    std_logic_vector(to_unsigned(192, n_bits_c)) when "11010100101", 
		    std_logic_vector(to_unsigned(193, n_bits_c)) when "11010100110", 
		    std_logic_vector(to_unsigned(194, n_bits_c)) when "11010100111", 
		    std_logic_vector(to_unsigned(195, n_bits_c)) when "11010101000", 
		    std_logic_vector(to_unsigned(196, n_bits_c)) when "11010101001", 
		    std_logic_vector(to_unsigned(197, n_bits_c)) when "11010101010", 
		    std_logic_vector(to_unsigned(197, n_bits_c)) when "11010101011", 
		    std_logic_vector(to_unsigned(198, n_bits_c)) when "11010101100", 
		    std_logic_vector(to_unsigned(199, n_bits_c)) when "11010101101", 
		    std_logic_vector(to_unsigned(200, n_bits_c)) when "11010101110", 
		    std_logic_vector(to_unsigned(201, n_bits_c)) when "11010101111", 
		    std_logic_vector(to_unsigned(202, n_bits_c)) when "11010110000", 
		    std_logic_vector(to_unsigned(202, n_bits_c)) when "11010110001", 
		    std_logic_vector(to_unsigned(203, n_bits_c)) when "11010110010", 
		    std_logic_vector(to_unsigned(204, n_bits_c)) when "11010110011", 
		    std_logic_vector(to_unsigned(205, n_bits_c)) when "11010110100", 
		    std_logic_vector(to_unsigned(206, n_bits_c)) when "11010110101", 
		    std_logic_vector(to_unsigned(207, n_bits_c)) when "11010110110", 
		    std_logic_vector(to_unsigned(208, n_bits_c)) when "11010110111", 
		    std_logic_vector(to_unsigned(209, n_bits_c)) when "11010111000", 
		    std_logic_vector(to_unsigned(210, n_bits_c)) when "11010111001", 
		    std_logic_vector(to_unsigned(210, n_bits_c)) when "11010111010", 
		    std_logic_vector(to_unsigned(211, n_bits_c)) when "11010111011", 
		    std_logic_vector(to_unsigned(212, n_bits_c)) when "11010111100", 
		    std_logic_vector(to_unsigned(213, n_bits_c)) when "11010111101", 
		    std_logic_vector(to_unsigned(214, n_bits_c)) when "11010111110", 
		    std_logic_vector(to_unsigned(215, n_bits_c)) when "11010111111", 
		    std_logic_vector(to_unsigned(216, n_bits_c)) when "11011000000", 
		    std_logic_vector(to_unsigned(217, n_bits_c)) when "11011000001", 
		    std_logic_vector(to_unsigned(218, n_bits_c)) when "11011000010", 
		    std_logic_vector(to_unsigned(219, n_bits_c)) when "11011000011", 
		    std_logic_vector(to_unsigned(220, n_bits_c)) when "11011000100", 
		    std_logic_vector(to_unsigned(221, n_bits_c)) when "11011000101", 
		    std_logic_vector(to_unsigned(222, n_bits_c)) when "11011000110", 
		    std_logic_vector(to_unsigned(222, n_bits_c)) when "11011000111", 
		    std_logic_vector(to_unsigned(223, n_bits_c)) when "11011001000", 
		    std_logic_vector(to_unsigned(224, n_bits_c)) when "11011001001", 
		    std_logic_vector(to_unsigned(225, n_bits_c)) when "11011001010", 
		    std_logic_vector(to_unsigned(226, n_bits_c)) when "11011001011", 
		    std_logic_vector(to_unsigned(227, n_bits_c)) when "11011001100", 
		    std_logic_vector(to_unsigned(228, n_bits_c)) when "11011001101", 
		    std_logic_vector(to_unsigned(229, n_bits_c)) when "11011001110", 
		    std_logic_vector(to_unsigned(230, n_bits_c)) when "11011001111", 
		    std_logic_vector(to_unsigned(231, n_bits_c)) when "11011010000", 
		    std_logic_vector(to_unsigned(232, n_bits_c)) when "11011010001", 
		    std_logic_vector(to_unsigned(233, n_bits_c)) when "11011010010", 
		    std_logic_vector(to_unsigned(234, n_bits_c)) when "11011010011", 
		    std_logic_vector(to_unsigned(235, n_bits_c)) when "11011010100", 
		    std_logic_vector(to_unsigned(236, n_bits_c)) when "11011010101", 
		    std_logic_vector(to_unsigned(237, n_bits_c)) when "11011010110", 
		    std_logic_vector(to_unsigned(238, n_bits_c)) when "11011010111", 
		    std_logic_vector(to_unsigned(239, n_bits_c)) when "11011011000", 
		    std_logic_vector(to_unsigned(240, n_bits_c)) when "11011011001", 
		    std_logic_vector(to_unsigned(241, n_bits_c)) when "11011011010", 
		    std_logic_vector(to_unsigned(242, n_bits_c)) when "11011011011", 
		    std_logic_vector(to_unsigned(243, n_bits_c)) when "11011011100", 
		    std_logic_vector(to_unsigned(244, n_bits_c)) when "11011011101", 
		    std_logic_vector(to_unsigned(246, n_bits_c)) when "11011011110", 
		    std_logic_vector(to_unsigned(247, n_bits_c)) when "11011011111", 
		    std_logic_vector(to_unsigned(248, n_bits_c)) when "11011100000", 
		    std_logic_vector(to_unsigned(249, n_bits_c)) when "11011100001", 
		    std_logic_vector(to_unsigned(250, n_bits_c)) when "11011100010", 
		    std_logic_vector(to_unsigned(251, n_bits_c)) when "11011100011", 
		    std_logic_vector(to_unsigned(252, n_bits_c)) when "11011100100", 
		    std_logic_vector(to_unsigned(253, n_bits_c)) when "11011100101", 
		    std_logic_vector(to_unsigned(254, n_bits_c)) when "11011100110", 
		    std_logic_vector(to_unsigned(255, n_bits_c)) when "11011100111", 
		    std_logic_vector(to_unsigned(256, n_bits_c)) when "11011101000", 
		    std_logic_vector(to_unsigned(257, n_bits_c)) when "11011101001", 
		    std_logic_vector(to_unsigned(258, n_bits_c)) when "11011101010", 
		    std_logic_vector(to_unsigned(260, n_bits_c)) when "11011101011", 
		    std_logic_vector(to_unsigned(261, n_bits_c)) when "11011101100", 
		    std_logic_vector(to_unsigned(262, n_bits_c)) when "11011101101", 
		    std_logic_vector(to_unsigned(263, n_bits_c)) when "11011101110", 
		    std_logic_vector(to_unsigned(264, n_bits_c)) when "11011101111", 
		    std_logic_vector(to_unsigned(265, n_bits_c)) when "11011110000", 
		    std_logic_vector(to_unsigned(266, n_bits_c)) when "11011110001", 
		    std_logic_vector(to_unsigned(267, n_bits_c)) when "11011110010", 
		    std_logic_vector(to_unsigned(268, n_bits_c)) when "11011110011", 
		    std_logic_vector(to_unsigned(270, n_bits_c)) when "11011110100", 
		    std_logic_vector(to_unsigned(271, n_bits_c)) when "11011110101", 
		    std_logic_vector(to_unsigned(272, n_bits_c)) when "11011110110", 
		    std_logic_vector(to_unsigned(273, n_bits_c)) when "11011110111", 
		    std_logic_vector(to_unsigned(274, n_bits_c)) when "11011111000", 
		    std_logic_vector(to_unsigned(275, n_bits_c)) when "11011111001", 
		    std_logic_vector(to_unsigned(276, n_bits_c)) when "11011111010", 
		    std_logic_vector(to_unsigned(278, n_bits_c)) when "11011111011", 
		    std_logic_vector(to_unsigned(279, n_bits_c)) when "11011111100", 
		    std_logic_vector(to_unsigned(280, n_bits_c)) when "11011111101", 
		    std_logic_vector(to_unsigned(281, n_bits_c)) when "11011111110", 
		    std_logic_vector(to_unsigned(282, n_bits_c)) when "11011111111", 
		    std_logic_vector(to_unsigned(283, n_bits_c)) when "11100000000", 
		    std_logic_vector(to_unsigned(285, n_bits_c)) when "11100000001", 
		    std_logic_vector(to_unsigned(286, n_bits_c)) when "11100000010", 
		    std_logic_vector(to_unsigned(287, n_bits_c)) when "11100000011", 
		    std_logic_vector(to_unsigned(288, n_bits_c)) when "11100000100", 
		    std_logic_vector(to_unsigned(289, n_bits_c)) when "11100000101", 
		    std_logic_vector(to_unsigned(291, n_bits_c)) when "11100000110", 
		    std_logic_vector(to_unsigned(292, n_bits_c)) when "11100000111", 
		    std_logic_vector(to_unsigned(293, n_bits_c)) when "11100001000", 
		    std_logic_vector(to_unsigned(294, n_bits_c)) when "11100001001", 
		    std_logic_vector(to_unsigned(295, n_bits_c)) when "11100001010", 
		    std_logic_vector(to_unsigned(297, n_bits_c)) when "11100001011", 
		    std_logic_vector(to_unsigned(298, n_bits_c)) when "11100001100", 
		    std_logic_vector(to_unsigned(299, n_bits_c)) when "11100001101", 
		    std_logic_vector(to_unsigned(300, n_bits_c)) when "11100001110", 
		    std_logic_vector(to_unsigned(302, n_bits_c)) when "11100001111", 
		    std_logic_vector(to_unsigned(303, n_bits_c)) when "11100010000", 
		    std_logic_vector(to_unsigned(304, n_bits_c)) when "11100010001", 
		    std_logic_vector(to_unsigned(305, n_bits_c)) when "11100010010", 
		    std_logic_vector(to_unsigned(306, n_bits_c)) when "11100010011", 
		    std_logic_vector(to_unsigned(308, n_bits_c)) when "11100010100", 
		    std_logic_vector(to_unsigned(309, n_bits_c)) when "11100010101", 
		    std_logic_vector(to_unsigned(310, n_bits_c)) when "11100010110", 
		    std_logic_vector(to_unsigned(311, n_bits_c)) when "11100010111", 
		    std_logic_vector(to_unsigned(313, n_bits_c)) when "11100011000", 
		    std_logic_vector(to_unsigned(314, n_bits_c)) when "11100011001", 
		    std_logic_vector(to_unsigned(315, n_bits_c)) when "11100011010", 
		    std_logic_vector(to_unsigned(317, n_bits_c)) when "11100011011", 
		    std_logic_vector(to_unsigned(318, n_bits_c)) when "11100011100", 
		    std_logic_vector(to_unsigned(319, n_bits_c)) when "11100011101", 
		    std_logic_vector(to_unsigned(320, n_bits_c)) when "11100011110", 
		    std_logic_vector(to_unsigned(322, n_bits_c)) when "11100011111", 
		    std_logic_vector(to_unsigned(323, n_bits_c)) when "11100100000", 
		    std_logic_vector(to_unsigned(324, n_bits_c)) when "11100100001", 
		    std_logic_vector(to_unsigned(326, n_bits_c)) when "11100100010", 
		    std_logic_vector(to_unsigned(327, n_bits_c)) when "11100100011", 
		    std_logic_vector(to_unsigned(328, n_bits_c)) when "11100100100", 
		    std_logic_vector(to_unsigned(329, n_bits_c)) when "11100100101", 
		    std_logic_vector(to_unsigned(331, n_bits_c)) when "11100100110", 
		    std_logic_vector(to_unsigned(332, n_bits_c)) when "11100100111", 
		    std_logic_vector(to_unsigned(333, n_bits_c)) when "11100101000", 
		    std_logic_vector(to_unsigned(335, n_bits_c)) when "11100101001", 
		    std_logic_vector(to_unsigned(336, n_bits_c)) when "11100101010", 
		    std_logic_vector(to_unsigned(337, n_bits_c)) when "11100101011", 
		    std_logic_vector(to_unsigned(339, n_bits_c)) when "11100101100", 
		    std_logic_vector(to_unsigned(340, n_bits_c)) when "11100101101", 
		    std_logic_vector(to_unsigned(341, n_bits_c)) when "11100101110", 
		    std_logic_vector(to_unsigned(343, n_bits_c)) when "11100101111", 
		    std_logic_vector(to_unsigned(344, n_bits_c)) when "11100110000", 
		    std_logic_vector(to_unsigned(345, n_bits_c)) when "11100110001", 
		    std_logic_vector(to_unsigned(347, n_bits_c)) when "11100110010", 
		    std_logic_vector(to_unsigned(348, n_bits_c)) when "11100110011", 
		    std_logic_vector(to_unsigned(349, n_bits_c)) when "11100110100", 
		    std_logic_vector(to_unsigned(351, n_bits_c)) when "11100110101", 
		    std_logic_vector(to_unsigned(352, n_bits_c)) when "11100110110", 
		    std_logic_vector(to_unsigned(353, n_bits_c)) when "11100110111", 
		    std_logic_vector(to_unsigned(355, n_bits_c)) when "11100111000", 
		    std_logic_vector(to_unsigned(356, n_bits_c)) when "11100111001", 
		    std_logic_vector(to_unsigned(357, n_bits_c)) when "11100111010", 
		    std_logic_vector(to_unsigned(359, n_bits_c)) when "11100111011", 
		    std_logic_vector(to_unsigned(360, n_bits_c)) when "11100111100", 
		    std_logic_vector(to_unsigned(362, n_bits_c)) when "11100111101", 
		    std_logic_vector(to_unsigned(363, n_bits_c)) when "11100111110", 
		    std_logic_vector(to_unsigned(364, n_bits_c)) when "11100111111", 
		    std_logic_vector(to_unsigned(366, n_bits_c)) when "11101000000", 
		    std_logic_vector(to_unsigned(367, n_bits_c)) when "11101000001", 
		    std_logic_vector(to_unsigned(369, n_bits_c)) when "11101000010", 
		    std_logic_vector(to_unsigned(370, n_bits_c)) when "11101000011", 
		    std_logic_vector(to_unsigned(371, n_bits_c)) when "11101000100", 
		    std_logic_vector(to_unsigned(373, n_bits_c)) when "11101000101", 
		    std_logic_vector(to_unsigned(374, n_bits_c)) when "11101000110", 
		    std_logic_vector(to_unsigned(376, n_bits_c)) when "11101000111", 
		    std_logic_vector(to_unsigned(377, n_bits_c)) when "11101001000", 
		    std_logic_vector(to_unsigned(378, n_bits_c)) when "11101001001", 
		    std_logic_vector(to_unsigned(380, n_bits_c)) when "11101001010", 
		    std_logic_vector(to_unsigned(381, n_bits_c)) when "11101001011", 
		    std_logic_vector(to_unsigned(383, n_bits_c)) when "11101001100", 
		    std_logic_vector(to_unsigned(384, n_bits_c)) when "11101001101", 
		    std_logic_vector(to_unsigned(385, n_bits_c)) when "11101001110", 
		    std_logic_vector(to_unsigned(387, n_bits_c)) when "11101001111", 
		    std_logic_vector(to_unsigned(388, n_bits_c)) when "11101010000", 
		    std_logic_vector(to_unsigned(390, n_bits_c)) when "11101010001", 
		    std_logic_vector(to_unsigned(391, n_bits_c)) when "11101010010", 
		    std_logic_vector(to_unsigned(393, n_bits_c)) when "11101010011", 
		    std_logic_vector(to_unsigned(394, n_bits_c)) when "11101010100", 
		    std_logic_vector(to_unsigned(395, n_bits_c)) when "11101010101", 
		    std_logic_vector(to_unsigned(397, n_bits_c)) when "11101010110", 
		    std_logic_vector(to_unsigned(398, n_bits_c)) when "11101010111", 
		    std_logic_vector(to_unsigned(400, n_bits_c)) when "11101011000", 
		    std_logic_vector(to_unsigned(401, n_bits_c)) when "11101011001", 
		    std_logic_vector(to_unsigned(403, n_bits_c)) when "11101011010", 
		    std_logic_vector(to_unsigned(404, n_bits_c)) when "11101011011", 
		    std_logic_vector(to_unsigned(406, n_bits_c)) when "11101011100", 
		    std_logic_vector(to_unsigned(407, n_bits_c)) when "11101011101", 
		    std_logic_vector(to_unsigned(409, n_bits_c)) when "11101011110", 
		    std_logic_vector(to_unsigned(410, n_bits_c)) when "11101011111", 
		    std_logic_vector(to_unsigned(411, n_bits_c)) when "11101100000", 
		    std_logic_vector(to_unsigned(413, n_bits_c)) when "11101100001", 
		    std_logic_vector(to_unsigned(414, n_bits_c)) when "11101100010", 
		    std_logic_vector(to_unsigned(416, n_bits_c)) when "11101100011", 
		    std_logic_vector(to_unsigned(417, n_bits_c)) when "11101100100", 
		    std_logic_vector(to_unsigned(419, n_bits_c)) when "11101100101", 
		    std_logic_vector(to_unsigned(420, n_bits_c)) when "11101100110", 
		    std_logic_vector(to_unsigned(422, n_bits_c)) when "11101100111", 
		    std_logic_vector(to_unsigned(423, n_bits_c)) when "11101101000", 
		    std_logic_vector(to_unsigned(425, n_bits_c)) when "11101101001", 
		    std_logic_vector(to_unsigned(426, n_bits_c)) when "11101101010", 
		    std_logic_vector(to_unsigned(428, n_bits_c)) when "11101101011", 
		    std_logic_vector(to_unsigned(429, n_bits_c)) when "11101101100", 
		    std_logic_vector(to_unsigned(431, n_bits_c)) when "11101101101", 
		    std_logic_vector(to_unsigned(432, n_bits_c)) when "11101101110", 
		    std_logic_vector(to_unsigned(434, n_bits_c)) when "11101101111", 
		    std_logic_vector(to_unsigned(435, n_bits_c)) when "11101110000", 
		    std_logic_vector(to_unsigned(437, n_bits_c)) when "11101110001", 
		    std_logic_vector(to_unsigned(438, n_bits_c)) when "11101110010", 
		    std_logic_vector(to_unsigned(440, n_bits_c)) when "11101110011", 
		    std_logic_vector(to_unsigned(441, n_bits_c)) when "11101110100", 
		    std_logic_vector(to_unsigned(443, n_bits_c)) when "11101110101", 
		    std_logic_vector(to_unsigned(444, n_bits_c)) when "11101110110", 
		    std_logic_vector(to_unsigned(446, n_bits_c)) when "11101110111", 
		    std_logic_vector(to_unsigned(447, n_bits_c)) when "11101111000", 
		    std_logic_vector(to_unsigned(449, n_bits_c)) when "11101111001", 
		    std_logic_vector(to_unsigned(450, n_bits_c)) when "11101111010", 
		    std_logic_vector(to_unsigned(452, n_bits_c)) when "11101111011", 
		    std_logic_vector(to_unsigned(454, n_bits_c)) when "11101111100", 
		    std_logic_vector(to_unsigned(455, n_bits_c)) when "11101111101", 
		    std_logic_vector(to_unsigned(457, n_bits_c)) when "11101111110", 
		    std_logic_vector(to_unsigned(458, n_bits_c)) when "11101111111", 
		    std_logic_vector(to_unsigned(460, n_bits_c)) when "11110000000", 
		    std_logic_vector(to_unsigned(461, n_bits_c)) when "11110000001", 
		    std_logic_vector(to_unsigned(463, n_bits_c)) when "11110000010", 
		    std_logic_vector(to_unsigned(464, n_bits_c)) when "11110000011", 
		    std_logic_vector(to_unsigned(466, n_bits_c)) when "11110000100", 
		    std_logic_vector(to_unsigned(467, n_bits_c)) when "11110000101", 
		    std_logic_vector(to_unsigned(469, n_bits_c)) when "11110000110", 
		    std_logic_vector(to_unsigned(470, n_bits_c)) when "11110000111", 
		    std_logic_vector(to_unsigned(472, n_bits_c)) when "11110001000", 
		    std_logic_vector(to_unsigned(474, n_bits_c)) when "11110001001", 
		    std_logic_vector(to_unsigned(475, n_bits_c)) when "11110001010", 
		    std_logic_vector(to_unsigned(477, n_bits_c)) when "11110001011", 
		    std_logic_vector(to_unsigned(478, n_bits_c)) when "11110001100", 
		    std_logic_vector(to_unsigned(480, n_bits_c)) when "11110001101", 
		    std_logic_vector(to_unsigned(481, n_bits_c)) when "11110001110", 
		    std_logic_vector(to_unsigned(483, n_bits_c)) when "11110001111", 
		    std_logic_vector(to_unsigned(485, n_bits_c)) when "11110010000", 
		    std_logic_vector(to_unsigned(486, n_bits_c)) when "11110010001", 
		    std_logic_vector(to_unsigned(488, n_bits_c)) when "11110010010", 
		    std_logic_vector(to_unsigned(489, n_bits_c)) when "11110010011", 
		    std_logic_vector(to_unsigned(491, n_bits_c)) when "11110010100", 
		    std_logic_vector(to_unsigned(492, n_bits_c)) when "11110010101", 
		    std_logic_vector(to_unsigned(494, n_bits_c)) when "11110010110", 
		    std_logic_vector(to_unsigned(496, n_bits_c)) when "11110010111", 
		    std_logic_vector(to_unsigned(497, n_bits_c)) when "11110011000", 
		    std_logic_vector(to_unsigned(499, n_bits_c)) when "11110011001", 
		    std_logic_vector(to_unsigned(500, n_bits_c)) when "11110011010", 
		    std_logic_vector(to_unsigned(502, n_bits_c)) when "11110011011", 
		    std_logic_vector(to_unsigned(503, n_bits_c)) when "11110011100", 
		    std_logic_vector(to_unsigned(505, n_bits_c)) when "11110011101", 
		    std_logic_vector(to_unsigned(507, n_bits_c)) when "11110011110", 
		    std_logic_vector(to_unsigned(508, n_bits_c)) when "11110011111", 
		    std_logic_vector(to_unsigned(510, n_bits_c)) when "11110100000", 
		    std_logic_vector(to_unsigned(511, n_bits_c)) when "11110100001", 
		    std_logic_vector(to_unsigned(513, n_bits_c)) when "11110100010", 
		    std_logic_vector(to_unsigned(515, n_bits_c)) when "11110100011", 
		    std_logic_vector(to_unsigned(516, n_bits_c)) when "11110100100", 
		    std_logic_vector(to_unsigned(518, n_bits_c)) when "11110100101", 
		    std_logic_vector(to_unsigned(519, n_bits_c)) when "11110100110", 
		    std_logic_vector(to_unsigned(521, n_bits_c)) when "11110100111", 
		    std_logic_vector(to_unsigned(523, n_bits_c)) when "11110101000", 
		    std_logic_vector(to_unsigned(524, n_bits_c)) when "11110101001", 
		    std_logic_vector(to_unsigned(526, n_bits_c)) when "11110101010", 
		    std_logic_vector(to_unsigned(527, n_bits_c)) when "11110101011", 
		    std_logic_vector(to_unsigned(529, n_bits_c)) when "11110101100", 
		    std_logic_vector(to_unsigned(531, n_bits_c)) when "11110101101", 
		    std_logic_vector(to_unsigned(532, n_bits_c)) when "11110101110", 
		    std_logic_vector(to_unsigned(534, n_bits_c)) when "11110101111", 
		    std_logic_vector(to_unsigned(536, n_bits_c)) when "11110110000", 
		    std_logic_vector(to_unsigned(537, n_bits_c)) when "11110110001", 
		    std_logic_vector(to_unsigned(539, n_bits_c)) when "11110110010", 
		    std_logic_vector(to_unsigned(540, n_bits_c)) when "11110110011", 
		    std_logic_vector(to_unsigned(542, n_bits_c)) when "11110110100", 
		    std_logic_vector(to_unsigned(544, n_bits_c)) when "11110110101", 
		    std_logic_vector(to_unsigned(545, n_bits_c)) when "11110110110", 
		    std_logic_vector(to_unsigned(547, n_bits_c)) when "11110110111", 
		    std_logic_vector(to_unsigned(548, n_bits_c)) when "11110111000", 
		    std_logic_vector(to_unsigned(550, n_bits_c)) when "11110111001", 
		    std_logic_vector(to_unsigned(552, n_bits_c)) when "11110111010", 
		    std_logic_vector(to_unsigned(553, n_bits_c)) when "11110111011", 
		    std_logic_vector(to_unsigned(555, n_bits_c)) when "11110111100", 
		    std_logic_vector(to_unsigned(557, n_bits_c)) when "11110111101", 
		    std_logic_vector(to_unsigned(558, n_bits_c)) when "11110111110", 
		    std_logic_vector(to_unsigned(560, n_bits_c)) when "11110111111", 
		    std_logic_vector(to_unsigned(562, n_bits_c)) when "11111000000", 
		    std_logic_vector(to_unsigned(563, n_bits_c)) when "11111000001", 
		    std_logic_vector(to_unsigned(565, n_bits_c)) when "11111000010", 
		    std_logic_vector(to_unsigned(566, n_bits_c)) when "11111000011", 
		    std_logic_vector(to_unsigned(568, n_bits_c)) when "11111000100", 
		    std_logic_vector(to_unsigned(570, n_bits_c)) when "11111000101", 
		    std_logic_vector(to_unsigned(571, n_bits_c)) when "11111000110", 
		    std_logic_vector(to_unsigned(573, n_bits_c)) when "11111000111", 
		    std_logic_vector(to_unsigned(575, n_bits_c)) when "11111001000", 
		    std_logic_vector(to_unsigned(576, n_bits_c)) when "11111001001", 
		    std_logic_vector(to_unsigned(578, n_bits_c)) when "11111001010", 
		    std_logic_vector(to_unsigned(580, n_bits_c)) when "11111001011", 
		    std_logic_vector(to_unsigned(581, n_bits_c)) when "11111001100", 
		    std_logic_vector(to_unsigned(583, n_bits_c)) when "11111001101", 
		    std_logic_vector(to_unsigned(585, n_bits_c)) when "11111001110", 
		    std_logic_vector(to_unsigned(586, n_bits_c)) when "11111001111", 
		    std_logic_vector(to_unsigned(588, n_bits_c)) when "11111010000", 
		    std_logic_vector(to_unsigned(589, n_bits_c)) when "11111010001", 
		    std_logic_vector(to_unsigned(591, n_bits_c)) when "11111010010", 
		    std_logic_vector(to_unsigned(593, n_bits_c)) when "11111010011", 
		    std_logic_vector(to_unsigned(594, n_bits_c)) when "11111010100", 
		    std_logic_vector(to_unsigned(596, n_bits_c)) when "11111010101", 
		    std_logic_vector(to_unsigned(598, n_bits_c)) when "11111010110", 
		    std_logic_vector(to_unsigned(599, n_bits_c)) when "11111010111", 
		    std_logic_vector(to_unsigned(601, n_bits_c)) when "11111011000", 
		    std_logic_vector(to_unsigned(603, n_bits_c)) when "11111011001", 
		    std_logic_vector(to_unsigned(604, n_bits_c)) when "11111011010", 
		    std_logic_vector(to_unsigned(606, n_bits_c)) when "11111011011", 
		    std_logic_vector(to_unsigned(608, n_bits_c)) when "11111011100", 
		    std_logic_vector(to_unsigned(609, n_bits_c)) when "11111011101", 
		    std_logic_vector(to_unsigned(611, n_bits_c)) when "11111011110", 
		    std_logic_vector(to_unsigned(613, n_bits_c)) when "11111011111", 
		    std_logic_vector(to_unsigned(614, n_bits_c)) when "11111100000", 
		    std_logic_vector(to_unsigned(616, n_bits_c)) when "11111100001", 
		    std_logic_vector(to_unsigned(618, n_bits_c)) when "11111100010", 
		    std_logic_vector(to_unsigned(619, n_bits_c)) when "11111100011", 
		    std_logic_vector(to_unsigned(621, n_bits_c)) when "11111100100", 
		    std_logic_vector(to_unsigned(623, n_bits_c)) when "11111100101", 
		    std_logic_vector(to_unsigned(624, n_bits_c)) when "11111100110", 
		    std_logic_vector(to_unsigned(626, n_bits_c)) when "11111100111", 
		    std_logic_vector(to_unsigned(628, n_bits_c)) when "11111101000", 
		    std_logic_vector(to_unsigned(629, n_bits_c)) when "11111101001", 
		    std_logic_vector(to_unsigned(631, n_bits_c)) when "11111101010", 
		    std_logic_vector(to_unsigned(633, n_bits_c)) when "11111101011", 
		    std_logic_vector(to_unsigned(634, n_bits_c)) when "11111101100", 
		    std_logic_vector(to_unsigned(636, n_bits_c)) when "11111101101", 
		    std_logic_vector(to_unsigned(638, n_bits_c)) when "11111101110", 
		    std_logic_vector(to_unsigned(639, n_bits_c)) when "11111101111", 
		    std_logic_vector(to_unsigned(641, n_bits_c)) when "11111110000", 
		    std_logic_vector(to_unsigned(643, n_bits_c)) when "11111110001", 
		    std_logic_vector(to_unsigned(644, n_bits_c)) when "11111110010", 
		    std_logic_vector(to_unsigned(646, n_bits_c)) when "11111110011", 
		    std_logic_vector(to_unsigned(648, n_bits_c)) when "11111110100", 
		    std_logic_vector(to_unsigned(649, n_bits_c)) when "11111110101", 
		    std_logic_vector(to_unsigned(651, n_bits_c)) when "11111110110", 
		    std_logic_vector(to_unsigned(653, n_bits_c)) when "11111110111", 
		    std_logic_vector(to_unsigned(654, n_bits_c)) when "11111111000", 
		    std_logic_vector(to_unsigned(656, n_bits_c)) when "11111111001", 
		    std_logic_vector(to_unsigned(658, n_bits_c)) when "11111111010", 
		    std_logic_vector(to_unsigned(659, n_bits_c)) when "11111111011", 
		    std_logic_vector(to_unsigned(661, n_bits_c)) when "11111111100", 
		    std_logic_vector(to_unsigned(663, n_bits_c)) when "11111111101", 
		    std_logic_vector(to_unsigned(664, n_bits_c)) when "11111111110", 
		    std_logic_vector(to_unsigned(666, n_bits_c)) when "11111111111", 
		    std_logic_vector(to_unsigned(667, n_bits_c)) when others;
    
end architecture tabela_sin;

